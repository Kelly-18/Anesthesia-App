��       �yellowbrick.regressor.residuals��ResidualsPlot���)��}�(�	is_fitted��auto��force_model���	estimator��sklearn.tree._classes��DecisionTreeRegressor���)��}�(�	criterion��squared_error��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K	�
n_outputs_�K�max_features_�K	�tree_��sklearn.tree._tree��Tree���K	�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h&�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C       �t�bK��R�}�(hK�
node_count�M��nodes�h%h(K ��h*��R�(KM���h/�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hDh2K ��hEh2K��hFh2K��hGh/�f8�����R�(Kh3NNNJ����J����K t�bK��hHhRK ��hIh2K(��hJhRK0��uK8KKt�b�Bj                           �F@�]����?           ��@       �                   �^@�Q��|�?D           @t@                          �Q@��+A�ȓ?�            �d@������������������������       �                     �?                          @Y@��XW7�?�            �d@                          �Q@ ���?             2@������������������������       �                     �?                          �D@ x?             1@	       
                 ��K@ ��W�h?             .@������������������������       �                     �?                          �C@  1f߻E?             ,@                          �R@      �<             *@������������������������       �                      @                        ��L@      �<             &@������������������������       �                     �?                          �S@      �<
             $@������������������������       �                     �?������������������������       �      ��	             "@������������������������       �      �<             �?                          �P@ &�G�zd?              @������������������������       �                     �?������������������������       �      ȼ             �?       2                    K@��p��?�            �b@                          �I@�����?             ?@                          �A@�"-���?             @������������������������       �                     @������������������������       �      м             @                          �O@ *\���x?             8@������������������������       �                     �?       +                   �S@ �Z�s?             7@       &                   �[@ T��6Z?             .@        #                   �V@ ����I?             (@!       "                   �Y@      �<
             $@������������������������       �                     �?������������������������       �      ��	             "@$       %                   @[@ (�G�zd?              @������������������������       �                     �?������������������������       �      ��             �?'       *                 03sJ@ ƚxV4b?             @(       )                 ��J@      �<              @������������������������       �                     �?������������������������       �                     �?������������������������       �      ��             �?,       /                   `U@ '��Q�~?              @-       .                   `[@      �<             @������������������������       �      �<             @������������������������       �      м              @0       1                     �?���xV4�?             @������������������������       �                      @������������������������       �      ��             �?3       J                   �M@�v��c��?u            @]@4       5                   �@@�r$<�6�?!            �@@������������������������       �                      @6       A                   @A@���O�m�?             9@7       8                    [@��p=
ד?              @������������������������       �                     @9       @                   �U@ ���Mb�?             @:       =                   @L@ ��Q�~?             @;       <                   �K@ �G�z�?              @������������������������       �                     �?������������������������       �      ��             �?>       ?                   @[@      �<              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �<             �?B       G                   `[@ �5�z}?             1@C       D                   `Y@ $-��t?             ,@������������������������       �                     �?E       F                   `T@ R�uhDg?             *@������������������������       �                     (@������������������������       �      �<             �?H       I                   �R@���xV4�?             @������������������������       �                     �?������������������������       �      ��              @K       X                    P@�~*:ǌ?T             U@L       O                   �Z@ >
ף�?             0@M       N                   �S@`�G�z�?             @������������������������       �                     �?������������������������       �      ��              @P       U                     �? @���ׄ?             *@Q       R                    �? ��xV4�?             @������������������������       �                     @S       T                 pfS@���xV4�?             @������������������������       �      ��              @������������������������       �                     �?V       W                   �[@ 8-��T?             @������������������������       �      ��             @������������������������       �      �<             �?Y       f                 pf�P@��aׁ?D             Q@Z       e                   �P@ U���q?             0@[       ^                    T@ p2�cd?             .@\       ]                   �R@  ��Q�~?             @������������������������       �      �<             @������������������������       �                     �?_       `                   �R@      �<             &@������������������������       �                     �?a       b                   �P@      �<
             $@������������������������       �      ��              @c       d                    Z@      �<              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �<             �?g       h                   `Z@ �R�ǡ�?4             J@������������������������       �                     @i       l                   �R@ |�j�?0             H@j       k                   @C@ ��xV4b?             @������������������������       �                     �?������������������������       �      ��              @m       �                    ]@ ��7�?-            �F@n       �                   �[@  �� �~?!            �@@o       ~                     �? � �G7|?             ?@p       u                   `Z@ ~
%#Z?             2@q       r                   `\@ ��xV4b?             @������������������������       �      ��             @s       t                    �?      �<              @������������������������       �                     �?������������������������       �                     �?v       {                    ?@ =L]n�?             (@w       z                   �S@ i�l�v?             @x       y                   �T@ ��xV4b?             @������������������������       �                      @������������������������       �                     �?������������������������       �      м             @|       }                   `P@ o�l�v?             @������������������������       �                     @������������������������       �      м             �?       �                   @E@ l�$%k?             *@�       �                    \@ ����I?             (@������������������������       �      ��	             "@�       �                   �Z@ ȚxV4b?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    \@      �<              @������������������������       �                     �?������������������������       �                     �?�       �                 @3�R@ a���}?             (@�       �                    A@  ��Q�~?              @������������������������       �                      @�       �                   �]@ l�l�v?             @������������������������       �                     @�       �                   @T@ ��xV4b?             @������������������������       �                      @������������������������       �      ��             �?������������������������       �                     @�       �                 03�L@ �= =~o?�            �c@�       �                    T@ fP@0 `?3            �I@�       �                    S@ *}���b?             &@������������������������       �                      @�       �                   `R@ ��jQ\?	             "@������������������������       �                     �?�       �                   �R@ P���Q?              @������������������������       �                     @�       �                   �V@ �G�zd?              @������������������������       �                     �?������������������������       �      ȼ             �?�       �                 ���L@ ,jM�S?(             D@�       �                    W@ Xx
E)N?'            �C@�       �                   �R@      �<             0@������������������������       �                     @�       �                   @V@      �<             &@������������������������       �                     �?������������������������       �      ȼ
             $@�       �                   @I@ �^�׉W?             7@������������������������       �                     �?�       �                    �? X��KS?             6@�       �                   pb@ �J�4a?
             $@�       �                   �V@  -��T?             @�       �                    W@ ��xV4b?             @������������������������       �                     �?������������������������       �      ��              @������������������������       �      ܼ             @�       �                    V@ ��xV4b?             @������������������������       �                     �?������������������������       �      ��              @�       �                   `W@      �<             (@������������������������       �                     @������������������������       �      ��             @������������������������       �                     �?�                         `V@ 8�I��n?j            �Z@�       �                 pf&M@ ��}�l?]            @W@�       �                   �V@ ��xV4b?             @������������������������       �                     �?�       �                   @S@      �<              @������������������������       �                     �?������������������������       �                     �?�       �                    �? �I��j?Z            �V@�       �                 `fS@ 贁Nk?0             H@�       �                 03�R@ �Qj�l?%            �B@�       �                   �V@ xffffd?              @@�       �                   �M@  ��Q�^?             0@�       �                     �? ��xV4b?             @������������������������       �      м              @������������������������       �      �<             �?�       �                 ��R@ x�k
TU?             *@������������������������       �      ��              @�       �                   `S@ @U0*�c?             @������������������������       �                      @�       �                   �a@ ��xV4b?             @������������������������       �                     �?������������������������       �      м              @�       �                   @U@ �����a?             0@�       �                   @C@ P���Q?              @������������������������       �                     @�       �                   @c@ �G�zd?              @������������������������       �                     �?������������������������       �      �<             �?�       �                    b@ �G�zd?              @������������������������       �                     @�       �                     �? 0��6Z?             @�       �                 ��9M@ �G�zd?              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �<             @�       �                    C@ �T0*�c?             @������������������������       �                      @�       �                   �R@      �<             @������������������������       �                     �?������������������������       �                      @�       �                 ��,T@ p�u_X?             &@�       �                    ?@ �H�}M?
             $@�       �                   �R@ �G�zd?              @������������������������       �                     �?������������������������       �                     �?������������������������       �      м              @������������������������       �                     �?�       �                   �U@ �&RN�g?*             E@������������������������       �                     @�       �                    R@ XD5X�e?'            �C@�       �                    W@ �G�zd?              @������������������������       �                     �?������������������������       �      ȼ             �?�       �                   �V@ h��c?%            �B@�       �                   @@@ �ZIfjY?             3@�       �                    b@ ��Q�^?              @�       �                   �a@      �<             @�       �                   �R@      �<              @������������������������       �                     �?������������������������       �                     �?������������������������       �      ��             �?�       �                   `V@ ,U0*�c?             @������������������������       �                      @�       �                   �W@      �<             @������������������������       �                     �?�       �                    ?@      �<              @������������������������       �                     �?������������������������       �                     �?�       �                 ���O@ ��߻K?             &@�       �                   �W@ ��xV4b?             @������������������������       �                     �?������������������������       �      ��              @������������������������       �      Լ              @�                       ��,Q@ ��0':d?             2@�                         �S@ h�l�V?             @�                          �V@ �G�zd?              @������������������������       �                     �?������������������������       �      �<             �?������������������������       �                     @                        �V@  ��Q�^?             (@������������������������       �                     �?      
                   V@ ��u_X?             &@                         S@ �H�}M?
             $@������������������������       �      м             @      	                  �S@ ��xV4b?             @������������������������       �                     �?������������������������       �      �<              @������������������������       �      �<             �?                        `b@ �uhDg?             *@������������������������       �                     @                        �W@ �H�}M?
             $@������������������������       �      ȼ	             "@������������������������       �                     �?      �                  `_@ \�^ŭ�?�             k@      G                   Q@ أ�`Έ?|             _@      F                `f�S@ ɐc�?2             I@      )                  �Z@ �S�ۇ?0             H@                         �? 
ᦛ?�?             7@                        @Y@ ~�Pk�?
             $@                        `X@ ��xV4b?             @������������������������       �                     �?������������������������       �                      @                        �S@ (-��t?             @������������������������       �                     @                        �Y@ �G�z�?              @������������������������       �                     �?������������������������       �      м             �?                         �N@ ��z�<x?             *@������������������������       �                     �?!      $                `f&N@ ؚxV4b?             (@"      #                  @K@ @��6Z?             @������������������������       �                     �?������������������������       �                     @%      &                ���N@      �<             @������������������������       �                     �?'      (                  �T@      �<             @������������������������       �                     �?������������������������       �                     @*      +                  @K@ �fh<�?             9@������������������������       �                     �?,      5                  �I@ �����z?             8@-      4                  @I@ (-��t?             @.      /                    �?      �<             @������������������������       �                     @0      1                  @W@      �<             @������������������������       �                     �?2      3                  �P@      �<              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �<             �?6      E                `f�R@ �����r?             1@7      <                  �K@ pffffn?             0@8      9                  �\@ `�l�V?             @������������������������       �                     @:      ;                   M@ �G�zd?              @������������������������       �                     �?������������������������       �      м             �?=      >                  `U@ �H�}m?
             $@������������������������       �                      @?      B                  �S@ �G�zd?              @@      A                  �P@ `�l�V?             @������������������������       �                     @������������������������       �      �<             �?C      D                    �? (�G�zd?              @������������������������       �                     �?������������������������       �      �<             �?������������������������       �      �             �?������������������������       �                      @H      O                `f&J@ ������?J            �R@I      L                  �Z@ �J�4a?
             $@J      K                  �X@  ��Q�^?             @������������������������       �                     �?������������������������       �                     @M      N                   S@      �<             @������������������������       �                     �?������������������������       �                     @P      c                  `R@ &��Q��?@             P@Q      b                  �W@ `�,{�?             9@R      _                   R@ lF!��?             7@S      T                  �R@ �_,�ł?             2@������������������������       �                      @U      \                   ]@ 23333�?             0@V      W                ��LM@ �h$��w?             (@������������������������       �                     @X      Y                  �H@ ���Mb�?             @������������������������       �                      @Z      [                  �V@ ��xV4b?             @������������������������       �                      @������������������������       �      �             �?]      ^                83�P@ 4��Q�~?             @������������������������       �      �             @������������������������       �                     �?`      a                    �?      �<             @������������������������       �                      @������������������������       �                     @������������������������       �      �              @d      �                  �Q@ J8�7��?'            �C@e      l                  @H@ |�j�?             8@f      g                  �P@ �G�z~?              @������������������������       �                     @h      i                ��iQ@ `���(|?             @������������������������       �                      @j      k                    �? �G�zd?              @������������������������       �                     �?������������������������       �      �<             �?m      �                  �]@  \���x?             0@n      o                  @K@ xT��r?             .@������������������������       �                     �?p      s                  �Y@ �0f߻e?             ,@q      r                    �? ��xV4�?             @������������������������       �                      @������������������������       �                     �?t      u                   P@      �<             &@������������������������       �                     �?v      w                  @L@      �<
             $@������������������������       �                     �?x      y                   U@      �<	             "@������������������������       �                     �?z      {                  �R@      �<              @������������������������       �                     �?|      }                `f�L@      �<             @������������������������       �                     �?~                        �Z@      �<             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                  �W@ Tn6��}?             .@�      �                  �H@ �%��`?             @������������������������       �                      @������������������������       �                     @�      �                   I@ f���(�?              @�      �                  �[@ �?^�k|?             @�      �                   S@ �G�z�?              @������������������������       �                     �?������������������������       �      м             �?�      �                  �S@ @��6Z?             @������������������������       �                     @������������������������       �      �             �?������������������������       �                     �?�      �                  `U@ ���|t?\             W@�      �                  �U@ �Ƞ7�q?S            �T@�      �                   R@ |�[V�q?#            �A@������������������������       �                      @�      �                    �? �S	 p?!            �@@�      �                  @L@ @^�kl?             ,@�      �                  @S@  -��T?             @������������������������       �      м             @������������������������       �                     �?�      �                ��lI@ �%��`?             @������������������������       �                     �?�      �                ���L@ @�l�V?             @�      �                03SL@ ��xV4b?             @������������������������       �                      @������������������������       �      �<             �?������������������������       �                     @�      �                  �P@ �r4�h?             3@�      �                  �R@ 贁Nk?             @�      �                  �R@  ��6Z?             @�      �                  �Q@ �G�zd?              @������������������������       �                     �?������������������������       �      �             �?�      �                  �N@      �<             @�      �                  �N@      �<              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �      �<             �?�      �                  �L@ �(b�cc?             *@�      �                  �R@ p��?`?             &@������������������������       �      м             @�      �                  `b@ HU0*�c?             @������������������������       �                      @������������������������       �      �             @������������������������       �       �              @�      �                  �R@ �����m?0             H@�      �                  �J@ �_�Le?(             D@�      �                  @J@ ����.p?	             "@�      �                    �? H3333c?              @�      �                  �R@ ��xV4b?             @������������������������       �                     �?������������������������       �                      @�      �                  `c@ `��6Z?             @������������������������       �                     �?������������������������       �                     @������������������������       �      �             �?�      �                  `S@ 0[Z�)V?             ?@�      �                  �c@ ����XO?             <@�      �                   S@ @��6Z?             .@�      �                  �R@ 03333c?              @������������������������       �                      @�      �                  �M@ p�l�V?             @������������������������       �                     @������������������������       �                     �?�      �                   �?      �<             @������������������������       �                     @������������������������       �      �             @�      �                   R@      �<             *@������������������������       �                     �?�      �                   �?      �<             (@������������������������       �      м              @�      �                  `R@      �<             @������������������������       �                     �?�      �                ��P@      �<             @�      �                  �c@      �<              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �                  �c@ H�xV4b?             @������������������������       �                      @������������������������       �      �             �?�      �                  `S@  \���x?              @������������������������       �                      @�      �                  �S@ �G�zd?             @�      �                  �c@      �<             @�      �                   T@      �<              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �      ��             @�      �                  @I@ آ�>7s?	             "@�      �                  �R@ ��xV4b?             @������������������������       �                     �?������������������������       �                      @�      �                   d@ ��l�V?             @������������������������       �                     @������������������������       �      ��             �?�t�b�values�h%h(K ��h*��R�(KM�KK��hR�B(  �e|���?q��g�?eK.�IE�?�������?x�G�5�?&}�'}��?ffffff�?233333�?�z�G��?      �?^�_��?233333�?333333�?233333�?333333�?233333�?333333�?333333�?�������?�������?�������?ffffff�?*�N��?���ۡ�?�_�_�?      �?333333�?�������?      �?���,d!�?��Q���?TUUUUU�?233333�?333333�?333333�?      �?333333�?�������?DDDDDD�?�������?�������?�������?333333�?ffffff�?333333�?333333�?333333�?�?      �?333333�?��؉���?߰�k��?      �?���x�&�?      �?      �?433333�?ffffff�?�������?333333�?      �?333333�?333333�?333333�?ffffff�?�������?PuPu�?333333�?�?�?�?      �?333333�?#"""""�?      �?333333�?��:��:�?������?gfffff�?�������?333333�?i�Vj�V�?�?      �?#"""""�?333333�?      �?۶m۶m�?333333�?�������?�?�������?�b�/���?ffffff�?333333�?      �?233333�?333333�?233333�?333333�?333333�?333333�?333333�?      �?��ȍ���?      �?�������?�������?�������?333333�?�i�6��?�[���?8z��'8�?q�q��?�������?333333�?�������?�������?�������?UUUUUU�?#"""""�?�?�������?      �?333333�?�������?      �?333333�?J��J���?�?333333�?�������?�������?333333�?      �?      �?      �?      �?�?�������?333333�?�?      �?#"""""�?�������?333333�?      �?=�T<׬�?�?b�־a�?ffffff�?}�'}�'�?ffffff�?      �?�������?�������?�������?ffffff�?D�z�G�?�c<�c<�?efffff�?ffffff�?gfffff�?ffffff�?gfffff�?aܯK*�?�������?,�袋.�?�Q����?��+��+�?�������?�������?ffffff�?ffffff�?UUUUUU�?ffffff�?�������?gfffff�?ffffff�?gfffff�?      �?�B�_��?�"�*�?�������?�������?      �?      �?      �?b�[��?333333�?�u�)�Y�?dffff&�?�������?xwwwww�?      �?ffffff�?Vj�Vj��?gfffff�?ףp=
�?ffffff�?xwwwww�?ffffff�?      �?     ��?�������?      �?333333�?      �?ffffff�?433333�?      �?���Q��?333333�?ffffff�?      �?efffff�?�p=
ף�?�������?      �?      �?      �?��k߰�?���(\��?333333�?ffffff�?      �?gfffff�?      �?�����?      �?�k��k��?�������?�������?ffffff�?��}M��?��8�{�?�������?efffff�?ffffff�?ffffff�?ffffff�?ffffff�?
ףp=
�?      �?efffff�?ffffff�?ffffff�?ffffff�?ffffff�?B��)A�?�������?�������?ffffff�?gfffff�?�q�q�?�������?333333�?      �?ffffff�?      �?�������?      �?��k߰�?���(\��?gfffff�?�������?      �?ffffff�?      �?vb'vb'�?�������?���(\��?gfffff�?      �?)j��#@@u;T�C@/�$�@�@V>��uI@���Q� @������@ffffff@������@��:��: @       @������ @       @������@����@       @������@=
ףp=@������@ffffff@������@������@������@������@������@m�����@       @gffff�@�_�_@������@������@������@������@������@������@������@       @@�����@������@������@      @������@ffffff@>
ףp=@������@ffffff@DDDDDD@ffffff@������@������@ffffff@333333@333333@       @�Qm�J@ףp=
�@333333@������@ffffff@������@������@������@������ @��S㥛 @�B��� @������ @������@����̌ @UUUUUU @       @������ @       @VUUUUU@������@������ @433333@������@       @       @       @       @������@�;�;@�����@     � @       @      @������@ffffff @������ @       @�����L@b�/��b@       @�W|�W|@@������@       @������@������@������@������@������@������@������@������@������@������@������@������@������@       @�%�X�@B�A�@ffffff@������@�����L@�W|�W|@������ @������@       @��(\��@������@ffffff@       @K[�#P@U�M�_@&�;Y-@ffffff@8��g9@������@uPuP@333333@      @��@333333@������@������@ffffff@333333@ffffff@�v�@i@333333@\���(\@������@333333@      @333333@333333@333333@333333@333333@ffffff@����@j߰�k@333333@�G�z�@333333@      @      @HDDDD�@s=
ףp@'}�'}�@33333�@wwwwww@      @333333@ףp=
�@333333@      @������@U�Cu;T@�$I�$I@[���(\@     �@      @UUUUUU@333333@      @333333@333333@333333@233333@333333@233333@333333@333333@333333@333333@333333@333333@333333@333333@������@      @333333@fffff�@������@������@333333@333333@333333@333333@333333@      @l�l�@""""""@������@ffffff@@333333@ffffff@�t�bub�_sklearn_version��1.0.2�ub�name�h
�_wrapped�h�_ax��matplotlib.axes._subplots��$_picklable_subplot_class_constructor����matplotlib.axes._axes��Axes�����R�}�(�_stale���stale_callback�N�_axes�hn�figure��matplotlib.figure��Figure���)��}�(hp�hqNhshw�
_transform�N�_transformSet���_visible���	_animated���_alpha�N�clipbox�N�	_clippath�N�_clipon���_label�� ��_picker�N�	_contains�N�_rasterized���_agg_filter�N�
_mouseover���
_callbacks��matplotlib.cbook��CallbackRegistry���)��}�(�exception_handler�h��_exception_printer����	callbacks�}��_cid_gen��	itertools��count���K ��R��_func_cid_map�N�_pickled_cids���ub�_remove_method�N�_url�N�_gid�N�_snap�N�_sketch�N�_path_effects�]��_sticky_edges��matplotlib.artist��_XYPair���]�]������
_in_layout���	_suptitle�N�
_supxlabel�N�
_supylabel�N�_align_label_groups�}�(�x�h��Grouper���)��}��_mapping�}�sb�y�h�)��}�h�}�sbu�
_gridspecs�]��
_localaxes�ht�
_AxesStack���)��}�(�_pos�K�	_elements�]�(Khn��Khl)��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh��builtins��getattr���hw�delaxes���R�h�Nh�Nh�Nh�Nh�h�h�h�]�]�����h���	_position��matplotlib.transforms��Bbox���)��}�(�_parents�}���]�hڌTransformedBbox���)��}�(h�}��]�hڌBboxTransformTo���)��}�(h�}�(��]�hڌCompositeGenericTransform���)��}�(�
input_dims�K�output_dims�Kh�}���]�h�)��}�(h�Kh�Kh�}�(� ]�hڌBlendedGenericTransform���)��}�(h�}�(�P^�h�)��}�(h�Kh�Kh�}��_invalid�K�_shorthand_name�h��_a�h��_b�hڌScaledTranslation���)��}�(h�}��P^�h�sh�K h�h��	_inverted�N�_t�K G���8�9���_scale_trans�hڌAffine2D���)��}�(h�}�(�0JM�h�)��}�(h�}���JM�h�)��}�(h�}�(� KW�h�)��}�(h�}����Z�h�)��}�(h�}�(���Z�h�)��}�(h�Kh�Kh�}����Z�h�)��}�(h�Kh�Kh�}�(���Z�h�)��}�(h�}�(���U�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j!  j   j  )��}�(h�}����U�j$  sh�K h�h�j  Nj  K G���8�9��j	  j  �_mtx�h%h(K ��h*��R�(KKK��hR�CH      �?                              �?      �                      �?�t�bubub���U�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j!  j   j  )��}�(h�}����U�j2  sh�Kh�h�j  Nj  K G?��8�9��j	  j  j+  Nubub���[�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j!  j   j  )��}�(h�}����[�j9  sh�K h�h�j  Nj  K G���8�9��j	  j  j+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?      �                      �?�t�bubub��[�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j!  j   j  )��}�(h�}���[�jF  sh�Kh�h�j  Nj  K G?��8�9��j	  j  j+  Nubub�0M\�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j!  j   j  )��}�(h�}��0M\�jM  sh�Kh�h�j  Nj  K G��-��-�؆�j	  j  j+  Nubub� J\�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j!  j   j  )��}�(h�}�� J\�jT  sh�Kh�h�j  Nj  K G?�-��-�؆�j	  j  j+  Nubub�`O�hڌTransformedPath���)��}�(h�}�h�Kh�h��_path��matplotlib.path��Path���)��}�(�	_vertices�h%h(K ��h*��R�(KKK��hR�C       �?      �?              �?�t�b�_codes�N�_interpolation_steps�K��_simplify_threshold�G?�q�q�֌_should_simplify���	_readonly��ubhyj!  �_transformed_path�jc  )��}�(jf  ji  jm  Njq  �jp  �jo  G?�q�q��jn  K�ub�_transformed_points�jc  )��}�(jf  ji  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub�PEM�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C 433333�?433333�?              �?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj!  jr  jc  )��}�(jf  j  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub���J�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C gfffff�?gfffff�?              �?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj!  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub�p�J�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C �������?�������?              �?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj!  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub��J�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C �������?�������?              �?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj!  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub�P�J�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C        @       @              �?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj!  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub�@`O�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C ������@������@              �?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj!  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub���J�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C 433333@433333@              �?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj!  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub��MM�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C ������@������@              �?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj!  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ububuh�Kh�h��_x�j  �_y�j  �_affine�j  )��}�(h�}�h�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CHt�E]�|@        �E]t�w�        ��(\�bt@������B@                      �?�t�bubub���Z�h�)��}�(h�}�(���[�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j�  j   j  )��}�(h�}����[�j�  sh�K h�h�j  Nj  G���8�9K ��j	  j  j+  h%h(K ��h*��R�(KKK��hR�CH      �?              �              �?                              �?�t�bubub�P�[�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j�  j   j  )��}�(h�}��P�[�j  sh�Kh�h�j  Nj  G?��8�9K ��j	  j  j+  Nubub��C\�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j�  j   j  )��}�(h�}���C\�j  sh�K h�h�j  Nj  G���8�9K ��j	  j  j+  h%h(K ��h*��R�(KKK��hR�CH      �?              �              �?                              �?�t�bubub��B\�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j�  j   j  )��}�(h�}���B\�j   sh�Kh�h�j  Nj  G?��8�9K ��j	  j  j+  Nubub��<\�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j�  j   j  )��}�(h�}���<\�j'  sh�Kh�h�j  Nj  G��-��-��K ��j	  j  j+  Nubub��6\�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j�  j   j  )��}�(h�}���6\�j.  sh�Kh�h�j  Nj  G?�-��-��K ��j	  j  j+  Nubub�p�M�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?                �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubhyj�  jr  jc  )��}�(jf  j<  jm  Njq  �jp  �jo  G?�q�q��jn  Kubju  jc  )��}�(jf  j<  jm  Njq  �jp  �jo  G?�q�q��jn  Kubub�/U�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?������ɿ������ɿ�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj�  jr  jc  )��}�(jf  jK  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  jK  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub� �J�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?                �t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj�  jr  jc  )��}�(jf  jZ  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  jZ  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub��;�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?�������?�������?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj�  jr  jc  )��}�(jf  ji  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  ji  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub�P�J�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?�������?�������?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj�  jr  jc  )��}�(jf  jx  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  jx  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub��-I�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?333333�?333333�?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyj�  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ububuh�Kh�h�j�  j  j�  j  j�  j  )��}�(h�}�h�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH�����l�@        �����	H@        ]t�E�t@:@���b@                      �?�t�bububuh�Kh�h�h�hڌTransformWrapper���)��}�(h�}�(���Z�h�)��}�(h�}����Z�hڌBboxTransformFrom���)��}�(h�}����Z�j  sh�K h�h�j  j  )��}�(h�}�h�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH*\���(�?        o=
ףp�?        �G�z��?�G�zֿ                      �?�t�bub�_boxin�j�  j+  h%h(K ��h*��R�(KKK��hR�CH.�袋.�?        �袋.��        �@�_)�?J6�d�M�?                      �?�t�bubsh�K h�h��_bbox�h�)��}�(h�}����Z�j�  sh�K h�h��_points�h%h(K ��h*��R�(KKK��hR�C p=
ףp�?�G�zֿq=
ףp@�p=
ף�?�t�b�_minpos�h%h(K ��h*��R�(KK��hR�C      �      ��t�b�_ignore���_points_orig�h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C p=
ףp�?�G�zֿq=
ףp@�p=
ף�?�t�bub���Z�j  uh�K h�h�h�Kh�K�_child�hڌBlendedAffine2D���)��}�(h�}����Z�j�  sh�K h�h�j�  hڌIdentityTransform���)��}�(h�}����X�j�  sh�Kh�h�j  Nubj�  j�  )��}�(h�}����X�j�  sh�Kh�h�j  Nubj  j  )��}�(h�}�h�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bub�	transform�h�j�  j�  ��R��transform_affine�h�j�  j�  ��R��transform_non_affine�h�j�  j�  ��R��transform_path�h�j�  j�  ��R��transform_path_affine�h�j�  j�  ��R��transform_path_non_affine�h�j�  j  ��R��
get_affine�h�j�  j  ��R��inverted�h�j�  j  ��R��
get_matrix�h�j�  j
  ��R�ubj   j  ubsh�Kh�h�h�j�  j   j  ub���Z�j!  ���Z�j�  ���Z�j�  )��}�(h�}�h�Kh�h�j�  j  j�  j�  )��}�(h�}����Z�j  sh�Kh�h�j  Nubj  Nj+  h%h(K ��h*��R�(KKK��hR�CH�����l�@        �����	H@              �?                              �?�t�bub�p�Z�j�  )��}�(h�}�h�Kh�h�j�  j  j�  j�  )��}�(h�}��p�Z�j  sh�Kh�h�j  Nubj  Nj+  h%h(K ��h*��R�(KKK��hR�CH�����l�@              b@              �?                              �?�t�bub�p�X�j�  )��}�(h�}�h�Kh�h�j�  j�  )��}�(h�}��p�X�j%  sh�Kh�h�j  Nubj�  j  j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                        ��(\�bt@������B@                      �?�t�bub�`�X�j�  )��}�(h�}�h�Kh�h�j�  j  j�  j�  )��}�(h�}��`�X�j1  sh�Kh�h�j  Nubj  Nj+  h%h(K ��h*��R�(KKK��hR�CH�����l�@              b@              �?                              �?�t�bub�@I\�h�)��}�(h�Kh�Kh�}��pI\�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��pI\�j@  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj=  j�  h%h(K ��h*��R�(KKK��hR�C       b@      K@������@��(\��w@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@I\�j=  sh�Kh�h�h�h�)��}�(h�}��I\�j^  sh�K h�h�j  N�_boxout�h�)��}�(h�}���H\�ja  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��I\�j^  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub�O\�h�)��}�(h�Kh�Kh�}��@O\�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��@O\�j�  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��O\�j�  sh�Kh�h�h�h�)��}�(h�}���N\�j�  sh�Kh�h�j  Njd  h�)��}�(h�}�� N\�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}���N\�j�  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub� �[�h�)��}�(h�Kh�Kh�}���0\�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���0\�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C �����	H@������B@gffff�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� �[�j�  sh�Kh�h�h�h�)��}�(h�}��0�[�j�  sh�K h�h�j  Njd  h�)��}�(h�}���O\�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��0�[�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub�`�Z�h�)��}�(h�Kh�Kh�}����Z�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����Z�j  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��`�Z�j  sh�Kh�h�h�h�)��}�(h�}��`j�j.  sh�Kh�h�j  Njd  h�)��}�(h�}��01\�j1  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}��`j�j.  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub��j�h�)��}�(h�Kh�Kh�}����K�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����K�jU  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjR  j�  h%h(K ��h*��R�(KKK��hR�C �����	H@������B@gffff�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���j�jR  sh�Kh�h�h�h�)��}�(h�}��Pj�js  sh�K h�h�j  Njd  h�)��}�(h�}��@�K�jv  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��Pj�js  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub�3\�h�)��}�(h�Kh�Kh�}��@3\�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��@3\�j�  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��3\�j�  sh�Kh�h�h�h�)��}�(h�}�� �:�j�  sh�Kh�h�j  Njd  h�)��}�(h�}���2\�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}�� �:�j�  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub��4\�h�)��}�(h�Kh�Kh�}���4\�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���4\�j�  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���4\�j�  sh�Kh�h�h�h�)��}�(h�}��`4\�j�  sh�Kh�h�j  Njd  h�)��}�(h�}���3\�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}��`4\�j�  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub��5\�h�)��}�(h�Kh�Kh�}��6\�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��6\�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj  j�  h%h(K ��h*��R�(KKK��hR�C       b@      K@������@��(\��w@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���5\�j  sh�Kh�h�h�h�)��}�(h�}���5\�j<  sh�K h�h�j  Njd  h�)��}�(h�}�� 5\�j?  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���5\�j<  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub�?\�h�)��}�(h�Kh�Kh�}��@?\�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��@?\�ji  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjf  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��?\�jf  sh�Kh�h�h�h�)��}�(h�}���>\�j�  sh�Kh�h�j  Njd  h�)��}�(h�}�� >\�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}���>\�j�  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub��]�h�)��}�(h�Kh�Kh�}�� ]�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� ]�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C �����	H@������B@gffff�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���]�j�  sh�Kh�h�h�h�)��}�(h�}���]�j�  sh�K h�h�j  Njd  h�)��}�(h�}���?\�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���]�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub�P]�h�)��}�(h�Kh�Kh�}���]�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���]�j�  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��P]�j�  sh�Kh�h�h�h�)��}�(h�}�� ]�j  sh�Kh�h�j  Njd  h�)��}�(h�}���]�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}�� ]�j  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub��]�h�)��}�(h�Kh�Kh�}�� ]�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� ]�j2  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj/  j�  h%h(K ��h*��R�(KKK��hR�C �����	H@������B@gffff�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���]�j/  sh�Kh�h�h�h�)��}�(h�}���]�jP  sh�K h�h�j  Njd  h�)��}�(h�}��]�jS  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���]�jP  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub�P]�h�)��}�(h�Kh�Kh�}���]�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���]�j}  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjz  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��P]�jz  sh�Kh�h�h�h�)��}�(h�}�� ]�j�  sh�Kh�h�j  Njd  h�)��}�(h�}���]�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}�� ]�j�  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub�9\�h�)��}�(h�Kh�Kh�}��@9\�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��@9\�j�  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��9\�j�  sh�Kh�h�h�h�)��}�(h�}���]�j�  sh�Kh�h�j  Njd  h�)��}�(h�}��]�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}���]�j�  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub�@c`�h�)��}�(h�Kh�Kh�}��pc`�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��pc`�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C �����	H@������B@gffff�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@c`�j�  sh�Kh�h�h�h�)��}�(h�}��c`�j  sh�K h�h�j  Njd  h�)��}�(h�}���b`�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��c`�j  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub��Of�h�)��}�(h�Kh�Kh�}���0��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���0��jF  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjC  j�  h%h(K ��h*��R�(KKK��hR�C �����	H@������B@gffff�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Of�jC  sh�Kh�h�h�h�)��}�(h�}���Of�jd  sh�K h�h�j  Njd  h�)��}�(h�}���Mf�jg  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���Of�jd  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ub�01��h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j  j   j  )��}�(h�}�(�01��j�  �0G\�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j  j   j�  ub�`G\�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�j  j   j�  ubuh�K h�h�j  Nj  G        G?�UUUUUU��j	  j  j+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?      @                      �?�t�bubub�0G\�j�  �`G\�j�  �p�M�h�)��}�(h�Kh�Kh�}��P�M�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��P�M�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C �����	H@������B@gffff�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��p�M�j�  sh�Kh�h�h�h�)��}�(h�}�� �M�j�  sh�K h�h�j  Njd  h�)��}�(h�}���N�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�� �M�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   j  ubuh�Kh�h�j  Njd  j  j+  h%h(K ��h*��R�(KKK��hR�CH�����l�@        �����	H@        ��(\�bt@������B@                      �?�t�bubsh�Kh�h�j�  h�)��}�(h�}�� KW�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C       �?      �?�������?)\���(�?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj  j�  h%h(K ��h*��R�(KKK��hR�C �����	H@������B@gffff�@�(\�µv@�t�bub��]�h�uh�Kh�h�j  Njd  j  j+  h%h(K ��h*��R�(KKK��hR�CH      �@        23333�W�              {@������0�                      �?�t�bubsh�K h�h�j�  h�)��}�(h�}��0JM�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       0@      @�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       0@      @�t�bubhyj  j�  h%h(K ��h*��R�(KKK��hR�C                       �@      {@�t�bub���X�j'  ���U�j5  �`�U�j<  ���[�jI  ��[�j  �м[�j  � �[�j  ��D\�j#  �P�U�jP  ��M\�jW  �0=\�j*  ��=\�j1  ���]�j  �^�j  )��}�(h�}��`^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�h�j   j.  ubsh�Kh�h�j  Nj  K G?��8�9��j	  j  j+  Nub��^�j  )��}�(h�}�� ^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�h�j   j5  ubsh�K h�h�j  Nj  K G���8�9��j	  j  j+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?      �                      �?�t�bub�p^�j  )��}�(h�}��@^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�h�j   jB  ubsh�Kh�h�j  Nj  K G?��8�9��j	  j  j+  Nub�@^�j  )��}�(h�}��p3^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�h�)��}�(h�}�(�p3^�jL  ��2^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�jO  j   j  )��}�(h�}���2^�jR  sh�K h�h�j  Nj  G?��8�9K ��j	  j  j+  h%h(K ��h*��R�(KKK��hR�CH      �?              @              �?                              �?�t�bubub�`:^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�jO  j   j  )��}�(h�}��`:^�j_  sh�Kh�h�j  Nj  G���8�9K ��j	  j  j+  Nubub�`4^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�jO  j   j  )��}�(h�}��`4^�jf  sh�K h�h�j  Nj  G?��8�9K ��j	  j  j+  h%h(K ��h*��R�(KKK��hR�CH      �?              @              �?                              �?�t�bubub�@�_�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�jO  j   j  )��}�(h�}��@�_�js  sh�Kh�h�j  Nj  G��-��-��K ��j	  j  j+  Nubub�p�_�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�jO  j   j  )��}�(h�}��p�_�jz  sh�Kh�h�j  Nj  G?�-��-��K ��j	  j  j+  Nubub���M�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?                �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubhyjO  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  Kubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  Kubub�01^�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?������ɿ������ɿ�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyjO  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub��J�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?                �t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyjO  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub� �H�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?�������?�������?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyjO  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub���I�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?�������?�������?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyjO  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubub��j�j\  )��}�(h�}�h�Kh�h�j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?333333�?333333�?�t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubhyjO  jr  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ubju  jc  )��}�(jf  j�  jm  Njq  �jp  �jo  G?�q�q��jn  K�ububuh�Kh�h�j�  h�j�  h�j�  j  )��}�(h�}�h�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH������Q@            '�@        ]t�E�t@:@���b@                      �?�t�bububj   jI  ubsh�Kh�h�j  Nj  G���8�9K ��j	  j  j+  Nub�04^�jU  ��:^�jb  ��;^�ji  �p<^�j  )��}�(h�}�(�P>^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�h�j   j�  ub��>^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�h�j   j�  ub��>^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�h�j   j�  ubuh�K h�h�j  Nj  G        G?�UUUUUU��j	  j  j+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?      @                      �?�t�bub���^�j  )��}�(h�}��`�^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�h�j   j�  ubsh�Kh�h�j  Nj  K G��-��-�؆�j	  j  j+  Nub���^�j  )��}�(h�}����^�h�)��}�(h�Kh�Kh�}�h�Kh�h�h�h�j   j�  ubsh�Kh�h�j  Nj  K G?�-��-�؆�j	  j  j+  Nub�Ц_�jv  ���_�j}  ��c`�j�  uh�K h�h�j  j  )��}�(h�}�h�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH�q�q�?                        �q�q�?                              �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      R@                              R@                              �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?      �                      �?�t�bubub�`^�j1  � ^�j8  �@^�jE  �`�^�j�  ���^�j	  uh�Kh�h�j�  h�j�  h�j�  j  )��}�(h�}�h�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH�$I�$I�?            '�@        ��(\�bt@������B@                      �?�t�bubub�0]�jO  uh�Kh�h�h�j�  )��}�(h�}�(��]�h�)��}�(h�}���]�j�  )��}�(h�}���]�h�sh�K h�h�j  j  )��}�(h�}�h�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH     �@                        �G�z��?�G�zֿ                      �?�t�bubj�  j'	  j+  h%h(K ��h*��R�(KKK��hR�CHAA`?               �        �@�_)�?J6�d�M�?                      �?�t�bubsh�K h�h�j�  h�)��}�(h�}���]�j'	  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C         �G�zֿ     �@�p=
ף�?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj$	  j�  h%h(K ��h*��R�(K�G      KK��hR�C         �G�zֿ     �@�p=
ף�?�t�bub��]�h�uh�K h�h�h�Kh�Kj�  j�  )��}�(h�}���]�j$	  sh�K h�h�j�  j�  )��}�(h�}�� �]�jW	  sh�Kh�h�j  Nubj�  j�  )��}�(h�}�� �]�jW	  sh�Kh�h�j  Nubj  j  )��}�(h�}�h�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj+  j�  ubj�  h�jW	  j�  ��R�j�  h�jW	  j�  ��R�j�  h�jW	  j�  ��R�j�  h�jW	  j�  ��R�j�  h�jW	  j�  ��R�j  h�jW	  j  ��R�j  h�jW	  j  ��R�j  h�jW	  j  ��R�j
  h�jW	  j
  ��R�ubj   h�ubsh�Kh�h�h�j*	  j   h�ub� ]�h��0]�jO  �`�]�j�  )��}�(h�}�h�Kh�h�j�  h�j�  j�  )��}�(h�}��`�]�j{	  sh�Kh�h�j  Nubj  Nj+  h%h(K ��h*��R�(KKK��hR�CH������Q@            '�@              �?                              �?�t�bub���]�j�  )��}�(h�}�h�Kh�h�j�  h�j�  j�  )��}�(h�}����]�j�	  sh�Kh�h�j  Nubj  Nj+  h%h(K ��h*��R�(KKK��hR�CH������Q@        gffff&�@              �?                              �?�t�bub� �]�j�  )��}�(h�}�h�Kh�h�j�  j�  )��}�(h�}�� �]�j�	  sh�Kh�h�j  Nubj�  h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                        ��(\�bt@      K@                      �?�t�bub�`�]�j�  )��}�(h�}�h�Kh�h�j�  h�j�  j�  )��}�(h�}��`�]�j�	  sh�Kh�h�j  Nubj  Nj+  h%h(K ��h*��R�(KKK��hR�CH������Q@        gffff&�@              �?                              �?�t�bub�P>^�j�  ��>^�j�  ��>^�j�  ���^�h�)��}�(h�Kh�Kh�}����^�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����^�j�	  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�	  j�  h%h(K ��h*��R�(KKK��hR�C gffff&�@      K@333333�@��(\��w@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����^�j�	  sh�Kh�h�h�h�)��}�(h�}��p�^�j�	  sh�K h�h�j  Njd  h�)��}�(h�}���?^�j�	  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��p�^�j�	  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���^�h�)��}�(h�Kh�Kh�}�� �^�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� �^�j�	  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�	  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����^�j�	  sh�Kh�h�h�h�)��}�(h�}����^�j
  sh�Kh�h�j  Njd  h�)��}�(h�}����^�j
  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}����^�j
  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� 7^�h�)��}�(h�Kh�Kh�}��07^�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��07^�j8
  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj5
  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� 7^�j5
  sh�Kh�h�h�h�)��}�(h�}���6^�jP
  sh�Kh�h�j  Njd  h�)��}�(h�}����^�jS
  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}���6^�jP
  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��^�h�)��}�(h�Kh�Kh�}�� ^�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� ^�jw
  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjt
  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���^�jt
  sh�Kh�h�h�h�)��}�(h�}��p^�j�
  sh�Kh�h�j  Njd  h�)��}�(h�}��6^�j�
  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}��p^�j�
  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��^�h�)��}�(h�Kh�Kh�}�� �^�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� �^�j�
  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�
  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���^�j�
  sh�Kh�h�h�h�)��}�(h�}����^�j�
  sh�Kh�h�j  Njd  h�)��}�(h�}�� �^�j�
  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}����^�j�
  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�p�^�h�)��}�(h�Kh�Kh�}����^�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����^�j�
  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�
  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��p�^�j�
  sh�Kh�h�h�h�)��}�(h�}��@�^�j  sh�Kh�h�j  Njd  h�)��}�(h�}����^�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}��@�^�j  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���^�h�)��}�(h�Kh�Kh�}�� �^�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� �^�j4  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj1  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����^�j1  sh�Kh�h�h�h�)��}�(h�}����^�jL  sh�Kh�h�j  Njd  h�)��}�(h�}��0�^�jO  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}����^�jL  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�@�^�h�)��}�(h�Kh�Kh�}��p�^�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��p�^�js  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjp  j�  h%h(K ��h*��R�(KKK��hR�C gffff&�@      K@333333�@��(\��w@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@�^�jp  sh�Kh�h�h�h�)��}�(h�}���^�j�  sh�K h�h�j  Njd  h�)��}�(h�}����^�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���^�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���_�h�)��}�(h�Kh�Kh�}���_�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���_�j�  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����_�j�  sh�Kh�h�h�h�)��}�(h�}����_�j�  sh�Kh�h�j  Njd  h�)��}�(h�}����_�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}����_�j�  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�0�_�h�)��}�(h�Kh�Kh�}��`�_�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��`�_�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��0�_�j�  sh�Kh�h�h�h�)��}�(h�}�� �_�j  sh�K h�h�j  Njd  h�)��}�(h�}��p�_�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�� �_�j  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���_�h�)��}�(h�Kh�Kh�}���_�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���_�jH  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjE  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����_�jE  sh�Kh�h�h�h�)��}�(h�}����_�j`  sh�Kh�h�j  Njd  h�)��}�(h�}���_�jc  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}����_�j`  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�0�_�h�)��}�(h�Kh�Kh�}��`�_�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��`�_�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��0�_�j�  sh�Kh�h�h�h�)��}�(h�}�� �_�j�  sh�K h�h�j  Njd  h�)��}�(h�}��p�_�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�� �_�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���_�h�)��}�(h�Kh�Kh�}���_�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���_�j�  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����_�j�  sh�Kh�h�h�h�)��}�(h�}����_�j�  sh�Kh�h�j  Njd  h�)��}�(h�}���_�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}����_�j�  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�p``�h�)��}�(h�Kh�Kh�}���``�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���``�j  sh�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj  j�  Nubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��p``�j  sh�Kh�h�h�h�)��}�(h�}��@``�j)  sh�Kh�h�j  Njd  h�)��}�(h�}��p�_�j,  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  Nubj   j  )��}�(h�}��@``�j)  sh�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�Ph`�h�)��}�(h�Kh�Kh�}���h`�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���h`�jP  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjM  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��Ph`�jM  sh�Kh�h�h�h�)��}�(h�}�� h`�jn  sh�K h�h�j  Njd  h�)��}�(h�}���g`�jq  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�� h`�jn  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��j`�h�)��}�(h�Kh�Kh�}���j`�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���j`�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���j`�j�  sh�Kh�h�h�h�)��}�(h�}���j`�j�  sh�K h�h�j  Njd  h�)��}�(h�}��i`�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���j`�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��l`�h�)��}�(h�Kh�Kh�}��l`�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��l`�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���l`�j�  sh�Kh�h�h�h�)��}�(h�}���l`�j  sh�K h�h�j  Njd  h�)��}�(h�}��Pk`�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���l`�j  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��n`�h�)��}�(h�Kh�Kh�}�� n`�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� n`�j1  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj.  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���n`�j.  sh�Kh�h�h�h�)��}�(h�}���n`�jO  sh�K h�h�j  Njd  h�)��}�(h�}��`m`�jR  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���n`�jO  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��`a�h�)��}�(h�Kh�Kh�}���`a�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���`a�j|  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjy  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���`a�jy  sh�Kh�h�h�h�)��}�(h�}��p`a�j�  sh�K h�h�j  Njd  h�)��}�(h�}��po`�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��p`a�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�@ca�h�)��}�(h�Kh�Kh�}���ba�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���ba�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@ca�j�  sh�Kh�h�h�h�)��}�(h�}��ca�j�  sh�K h�h�j  Njd  h�)��}�(h�}���aa�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��ca�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�Pea�h�)��}�(h�Kh�Kh�}���da�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���da�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��Pea�j  sh�Kh�h�h�h�)��}�(h�}�� ea�j0  sh�K h�h�j  Njd  h�)��}�(h�}���ca�j3  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�� ea�j0  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�`ga�h�)��}�(h�Kh�Kh�}���fa�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���fa�j]  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjZ  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��`ga�jZ  sh�Kh�h�h�h�)��}�(h�}��0ga�j{  sh�K h�h�j  Njd  h�)��}�(h�}���ea�j~  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��0ga�j{  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��ha�h�)��}�(h�Kh�Kh�}���ha�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���ha�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���ha�j�  sh�Kh�h�h�h�)��}�(h�}���ga�j�  sh�K h�h�j  Njd  h�)��}�(h�}���ga�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���ga�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��ja�h�)��}�(h�Kh�Kh�}��0ja�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��0ja�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���ja�j�  sh�Kh�h�h�h�)��}�(h�}���ja�j  sh�K h�h�j  Njd  h�)��}�(h�}��pia�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���ja�j  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� ma�h�)��}�(h�Kh�Kh�}��@la�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��@la�j>  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj;  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� ma�j;  sh�Kh�h�h�h�)��}�(h�}���la�j\  sh�K h�h�j  Njd  h�)��}�(h�}���ka�j_  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���la�j\  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�oa�h�)��}�(h�Kh�Kh�}��Pna�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��Pna�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��oa�j�  sh�Kh�h�h�h�)��}�(h�}���na�j�  sh�K h�h�j  Njd  h�)��}�(h�}���ma�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���na�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��pb�h�)��}�(h�Kh�Kh�}�� qb�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� qb�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���pb�j�  sh�Kh�h�h�h�)��}�(h�}���pb�j�  sh�K h�h�j  Njd  h�)��}�(h�}���oa�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���pb�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�psb�h�)��}�(h�Kh�Kh�}���rb�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���rb�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��psb�j  sh�Kh�h�h�h�)��}�(h�}��@sb�j=  sh�K h�h�j  Njd  h�)��}�(h�}���qb�j@  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��@sb�j=  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��ub�h�)��}�(h�Kh�Kh�}���tb�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���tb�jj  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjg  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���ub�jg  sh�Kh�h�h�h�)��}�(h�}��Pub�j�  sh�K h�h�j  Njd  h�)��}�(h�}�� tb�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��Pub�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��wb�h�)��}�(h�Kh�Kh�}���vb�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���vb�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���wb�j�  sh�Kh�h�h�h�)��}�(h�}��`wb�j�  sh�K h�h�j  Njd  h�)��}�(h�}��vb�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��`wb�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��yb�h�)��}�(h�Kh�Kh�}���xb�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���xb�j   sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���yb�j�  sh�Kh�h�h�h�)��}�(h�}��pyb�j  sh�K h�h�j  Njd  h�)��}�(h�}�� xb�j!  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��pyb�j  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��{b�h�)��}�(h�Kh�Kh�}���zb�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���zb�jK  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjH  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���{b�jH  sh�Kh�h�h�h�)��}�(h�}���{b�ji  sh�K h�h�j  Njd  h�)��}�(h�}��0zb�jl  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���{b�ji  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��}b�h�)��}�(h�Kh�Kh�}�� }b�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� }b�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���}b�j�  sh�Kh�h�h�h�)��}�(h�}���}b�j�  sh�K h�h�j  Njd  h�)��}�(h�}��@|b�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���}b�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��b�h�)��}�(h�Kh�Kh�}��b�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��b�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���b�j�  sh�Kh�h�h�h�)��}�(h�}���b�j�  sh�K h�h�j  Njd  h�)��}�(h�}��P~b�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���b�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� Rc�h�)��}�(h�Kh�Kh�}��`Qc�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��`Qc�j,  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj)  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� Rc�j)  sh�Kh�h�h�h�)��}�(h�}���Qc�jJ  sh�K h�h�j  Njd  h�)��}�(h�}��@Pc�jM  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���Qc�jJ  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�0Tc�h�)��}�(h�Kh�Kh�}��pSc�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��pSc�jw  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjt  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��0Tc�jt  sh�Kh�h�h�h�)��}�(h�}�� Tc�j�  sh�K h�h�j  Njd  h�)��}�(h�}���Rc�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�� Tc�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�@Vc�h�)��}�(h�Kh�Kh�}���Uc�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Uc�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@Vc�j�  sh�Kh�h�h�h�)��}�(h�}��Vc�j�  sh�K h�h�j  Njd  h�)��}�(h�}���Tc�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��Vc�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�PXc�h�)��}�(h�Kh�Kh�}���Wc�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Wc�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj
  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��PXc�j
  sh�Kh�h�h�h�)��}�(h�}�� Xc�j+  sh�K h�h�j  Njd  h�)��}�(h�}���Vc�j.  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�� Xc�j+  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�`Zc�h�)��}�(h�Kh�Kh�}���Yc�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Yc�jX  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjU  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��`Zc�jU  sh�Kh�h�h�h�)��}�(h�}��0Zc�jv  sh�K h�h�j  Njd  h�)��}�(h�}���Xc�jy  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��0Zc�jv  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�p\c�h�)��}�(h�Kh�Kh�}���[c�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���[c�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��p\c�j�  sh�Kh�h�h�h�)��}�(h�}��@\c�j�  sh�K h�h�j  Njd  h�)��}�(h�}���Zc�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��@\c�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��^c�h�)��}�(h�Kh�Kh�}���]c�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���]c�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���^c�j�  sh�Kh�h�h�h�)��}�(h�}��P^c�j  sh�K h�h�j  Njd  h�)��}�(h�}�� ]c�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��P^c�j  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��`d�h�)��}�(h�Kh�Kh�}��p`d�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��p`d�j9  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj6  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���`d�j6  sh�Kh�h�h�h�)��}�(h�}��p_c�jW  sh�K h�h�j  Njd  h�)��}�(h�}��_c�jZ  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��p_c�jW  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��bd�h�)��}�(h�Kh�Kh�}�� bd�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� bd�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���bd�j�  sh�Kh�h�h�h�)��}�(h�}���bd�j�  sh�K h�h�j  Njd  h�)��}�(h�}��`ad�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���bd�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��dd�h�)��}�(h�Kh�Kh�}��0dd�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��0dd�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���dd�j�  sh�Kh�h�h�h�)��}�(h�}���dd�j�  sh�K h�h�j  Njd  h�)��}�(h�}��pcd�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���dd�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� gd�h�)��}�(h�Kh�Kh�}��@fd�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��@fd�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� gd�j  sh�Kh�h�h�h�)��}�(h�}���fd�j8  sh�K h�h�j  Njd  h�)��}�(h�}���ed�j;  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���fd�j8  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�id�h�)��}�(h�Kh�Kh�}��Phd�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��Phd�je  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjb  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��id�jb  sh�Kh�h�h�h�)��}�(h�}���hd�j�  sh�K h�h�j  Njd  h�)��}�(h�}���gd�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���hd�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� kd�h�)��}�(h�Kh�Kh�}��`jd�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��`jd�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� kd�j�  sh�Kh�h�h�h�)��}�(h�}���jd�j�  sh�K h�h�j  Njd  h�)��}�(h�}���id�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���jd�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�0md�h�)��}�(h�Kh�Kh�}��pld�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��pld�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��0md�j�  sh�Kh�h�h�h�)��}�(h�}�� md�j  sh�K h�h�j  Njd  h�)��}�(h�}���kd�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�� md�j  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�@od�h�)��}�(h�Kh�Kh�}���nd�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���nd�jF  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjC  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@od�jC  sh�Kh�h�h�h�)��}�(h�}��od�jd  sh�K h�h�j  Njd  h�)��}�(h�}���md�jg  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��od�jd  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Ae�h�)��}�(h�Kh�Kh�}���@e�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���@e�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Ae�j�  sh�Kh�h�h�h�)��}�(h�}��`Ae�j�  sh�K h�h�j  Njd  h�)��}�(h�}��@@e�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��`Ae�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Ce�h�)��}�(h�Kh�Kh�}���Be�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Be�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Ce�j�  sh�Kh�h�h�h�)��}�(h�}��pCe�j�  sh�K h�h�j  Njd  h�)��}�(h�}�� Be�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��pCe�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Ee�h�)��}�(h�Kh�Kh�}���De�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���De�j'  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj$  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Ee�j$  sh�Kh�h�h�h�)��}�(h�}���Ee�jE  sh�K h�h�j  Njd  h�)��}�(h�}��0De�jH  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���Ee�jE  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Ge�h�)��}�(h�Kh�Kh�}�� Ge�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� Ge�jr  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjo  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Ge�jo  sh�Kh�h�h�h�)��}�(h�}���Ge�j�  sh�K h�h�j  Njd  h�)��}�(h�}��@Fe�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���Ge�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Ie�h�)��}�(h�Kh�Kh�}��Ie�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��Ie�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Ie�j�  sh�Kh�h�h�h�)��}�(h�}���Ie�j�  sh�K h�h�j  Njd  h�)��}�(h�}��PHe�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���Ie�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Ke�h�)��}�(h�Kh�Kh�}�� Ke�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� Ke�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Ke�j  sh�Kh�h�h�h�)��}�(h�}���Ke�j&  sh�K h�h�j  Njd  h�)��}�(h�}��`Je�j)  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���Ke�j&  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Me�h�)��}�(h�Kh�Kh�}��0Me�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��0Me�jS  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjP  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Me�jP  sh�Kh�h�h�h�)��}�(h�}���Me�jq  sh�K h�h�j  Njd  h�)��}�(h�}��pLe�jt  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���Me�jq  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�@Oe�h�)��}�(h�Kh�Kh�}���Ne�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Ne�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@Oe�j�  sh�Kh�h�h�h�)��}�(h�}���Oe�j�  sh�K h�h�j  Njd  h�)��}�(h�}���Ne�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���Oe�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Af�h�)��}�(h�Kh�Kh�}���Af�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Af�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Af�j�  sh�Kh�h�h�h�)��}�(h�}���Af�j  sh�K h�h�j  Njd  h�)��}�(h�}�� Af�j
  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���Af�j  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�`Df�h�)��}�(h�Kh�Kh�}���Cf�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Cf�j4  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj1  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��`Df�j1  sh�Kh�h�h�h�)��}�(h�}��0Df�jR  sh�K h�h�j  Njd  h�)��}�(h�}���Bf�jU  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��0Df�jR  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�pFf�h�)��}�(h�Kh�Kh�}���Ef�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Ef�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj|  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��pFf�j|  sh�Kh�h�h�h�)��}�(h�}��@Ff�j�  sh�K h�h�j  Njd  h�)��}�(h�}���Df�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��@Ff�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Hf�h�)��}�(h�Kh�Kh�}���Gf�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Gf�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Hf�j�  sh�Kh�h�h�h�)��}�(h�}��PHf�j�  sh�K h�h�j  Njd  h�)��}�(h�}�� Gf�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��PHf�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Jf�h�)��}�(h�Kh�Kh�}���If�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���If�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Jf�j  sh�Kh�h�h�h�)��}�(h�}��`Jf�j3  sh�K h�h�j  Njd  h�)��}�(h�}��If�j6  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��`Jf�j3  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Lf�h�)��}�(h�Kh�Kh�}���Kf�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Kf�j`  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj]  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Lf�j]  sh�Kh�h�h�h�)��}�(h�}��pLf�j~  sh�K h�h�j  Njd  h�)��}�(h�}�� Kf�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��pLf�j~  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��Nf�h�)��}�(h�Kh�Kh�}���Mf�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���Mf�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���Nf�j�  sh�Kh�h�h�h�)��}�(h�}���Nf�j�  sh�K h�h�j  Njd  h�)��}�(h�}��0Mf�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���Nf�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� 5��h�)��}�(h�Kh�Kh�}��P5��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��P5��j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� 5��j�  sh�Kh�h�h�h�)��}�(h�}���4��j  sh�K h�h�j  Njd  h�)��}�(h�}��`4��j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���4��j  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��7��h�)��}�(h�Kh�Kh�}���7��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���7��jA  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj>  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���7��j>  sh�Kh�h�h�h�)��}�(h�}��`7��j_  sh�K h�h�j  Njd  h�)��}�(h�}���5��jb  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��`7��j_  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��9��h�)��}�(h�Kh�Kh�}���8��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���8��j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���9��j�  sh�Kh�h�h�h�)��}�(h�}��p9��j�  sh�K h�h�j  Njd  h�)��}�(h�}�� 8��j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��p9��j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubub�	      j   h�ub��;��h�)��}�(h�Kh�Kh�}���:��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���:��j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���;��j�  sh�Kh�h�h�h�)��}�(h�}���;��j�  sh�K h�h�j  Njd  h�)��}�(h�}��0:��j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���;��j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��=��h�)��}�(h�Kh�Kh�}�� =��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� =��j"  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���=��j  sh�Kh�h�h�h�)��}�(h�}���=��j@  sh�K h�h�j  Njd  h�)��}�(h�}��@<��jC  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���=��j@  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��?��h�)��}�(h�Kh�Kh�}��?��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��?��jm  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjj  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���?��jj  sh�Kh�h�h�h�)��}�(h�}���?��j�  sh�K h�h�j  Njd  h�)��}�(h�}��P>��j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���?��j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub����h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�����j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�����j�  sh�Kh�h�h�h�)��}�(h�}��`��j�  sh�K h�h�j  Njd  h�)��}�(h�}��� ��j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��`��j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�0��h�)��}�(h�Kh�Kh�}��p��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��p��j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj   j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��0��j   sh�Kh�h�h�h�)��}�(h�}�� ��j!  sh�K h�h�j  Njd  h�)��}�(h�}�����j$  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�� ��j!  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�@��h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�����jN  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjK  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@��jK  sh�Kh�h�h�h�)��}�(h�}����jl  sh�K h�h�j  Njd  h�)��}�(h�}�����jo  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}����jl  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�PK\�h�)��}�(h�Kh�Kh�}���L\�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���L\�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��PK\�j�  sh�Kh�h�h�h�)��}�(h�}���^�j�  sh�K h�h�j  Njd  h�)��}�(h�}���^�j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���^�j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���X�h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�����j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����X�j�  sh�Kh�h�h�h�)��}�(h�}��p�X�j  sh�K h�h�j  Njd  h�)��}�(h�}����X�j  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��p�X�j  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub����h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�����j/  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj,  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�����j,  sh�Kh�h�h�h�)��}�(h�}��P��jM  sh�K h�h�j  Njd  h�)��}�(h�}�� ��jP  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��P��jM  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��
��h�)��}�(h�Kh�Kh�}���	��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���	��jz  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjw  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���
��jw  sh�Kh�h�h�h�)��}�(h�}��`
��j�  sh�K h�h�j  Njd  h�)��}�(h�}��	��j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��`
��j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub����h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�����j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�����j�  sh�Kh�h�h�h�)��}�(h�}��p��j�  sh�K h�h�j  Njd  h�)��}�(h�}�� ��j�  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��p��j�  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub����h�)��}�(h�Kh�Kh�}�����h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�����j   sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj   j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�����j   sh�Kh�h�h�h�)��}�(h�}�����j.   sh�K h�h�j  Njd  h�)��}�(h�}��0��j1   sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�����j.   sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�p0��h�)��}�(h�Kh�Kh�}���0��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���0��j[   sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjX   j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��p0��jX   sh�Kh�h�h�h�)��}�(h�}��@0��jy   sh�K h�h�j  Njd  h�)��}�(h�}��@��j|   sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��@0��jy   sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�3��h�)��}�(h�Kh�Kh�}��P2��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��P2��j�   sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�   j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��3��j�   sh�Kh�h�h�h�)��}�(h�}���2��j�   sh�K h�h�j  Njd  h�)��}�(h�}���1��j�   sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���2��j�   sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� 5��h�)��}�(h�Kh�Kh�}��`4��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��`4��j�   sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�   j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� 5��j�   sh�Kh�h�h�h�)��}�(h�}���4��j!  sh�K h�h�j  Njd  h�)��}�(h�}���3��j!  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���4��j!  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�07��h�)��}�(h�Kh�Kh�}��p6��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��p6��j<!  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj9!  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��07��j9!  sh�Kh�h�h�h�)��}�(h�}�� 7��jZ!  sh�K h�h�j  Njd  h�)��}�(h�}���5��j]!  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}�� 7��jZ!  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�@9��h�)��}�(h�Kh�Kh�}���8��h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���8��j�!  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�!  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@9��j�!  sh�Kh�h�h�h�)��}�(h�}��9��j�!  sh�K h�h�j  Njd  h�)��}�(h�}���7��j�!  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��9��j�!  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�P�V�h�)��}�(h�Kh�Kh�}��@�W�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��@�W�j�!  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�!  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��P�V�j�!  sh�Kh�h�h�h�)��}�(h�}����V�j�!  sh�K h�h�j  Njd  h�)��}�(h�}����V�j�!  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}����V�j�!  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���X�h�)��}�(h�Kh�Kh�}��P�X�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��P�X�j"  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj"  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����X�j"  sh�Kh�h�h�h�)��}�(h�}��@�W�j;"  sh�K h�h�j  Njd  h�)��}�(h�}��p�W�j>"  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��@�W�j;"  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�P�X�h�)��}�(h�Kh�Kh�}����X�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����X�jh"  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyje"  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��P�X�je"  sh�Kh�h�h�h�)��}�(h�}��P�X�j�"  sh�K h�h�j  Njd  h�)��}�(h�}���X�j�"  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��P�X�j�"  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� �X�h�)��}�(h�Kh�Kh�}����X�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����X�j�"  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�"  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� �X�j�"  sh�Kh�h�h�h�)��}�(h�}����X�j�"  sh�K h�h�j  Njd  h�)��}�(h�}���X�j�"  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}����X�j�"  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�0�W�h�)��}�(h�Kh�Kh�}���W�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���W�j�"  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�"  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��0�W�j�"  sh�Kh�h�h�h�)��}�(h�}��@�W�j#  sh�K h�h�j  Njd  h�)��}�(h�}����W�j#  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��@�W�j#  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���W�h�)��}�(h�Kh�Kh�}���W�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���W�jI#  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjF#  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����W�jF#  sh�Kh�h�h�h�)��}�(h�}����W�jg#  sh�K h�h�j  Njd  h�)��}�(h�}��`�W�jj#  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}����W�jg#  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�pCW�h�)��}�(h�Kh�Kh�}��@FW�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��@FW�j�#  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�#  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��pCW�j�#  sh�Kh�h�h�h�)��}�(h�}��@CW�j�#  sh�K h�h�j  Njd  h�)��}�(h�}���NW�j�#  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��@CW�j�#  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� �T�h�)��}�(h�Kh�Kh�}��@�T�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��@�T�j�#  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�#  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� �T�j�#  sh�Kh�h�h�h�)��}�(h�}����T�j�#  sh�K h�h�j  Njd  h�)��}�(h�}��OW�j $  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}����T�j�#  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�P�T�h�)��}�(h�Kh�Kh�}��МT�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��МT�j*$  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj'$  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��P�T�j'$  sh�Kh�h�h�h�)��}�(h�}����T�jH$  sh�K h�h�j  Njd  h�)��}�(h�}��0�T�jK$  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}����T�jH$  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���K�h�)��}�(h�Kh�Kh�}�� �K�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� �K�ju$  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjr$  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����K�jr$  sh�Kh�h�h�h�)��}�(h�}��0�K�j�$  sh�K h�h�j  Njd  h�)��}�(h�}����K�j�$  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��0�K�j�$  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���K�h�)��}�(h�Kh�Kh�}����K�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����K�j�$  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�$  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����K�j�$  sh�Kh�h�h�h�)��}�(h�}��`�K�j�$  sh�K h�h�j  Njd  h�)��}�(h�}����K�j�$  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��`�K�j�$  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�@�K�h�)��}�(h�Kh�Kh�}��p�K�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��p�K�j%  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj%  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@�K�j%  sh�Kh�h�h�h�)��}�(h�}��0�K�j)%  sh�K h�h�j  Njd  h�)��}�(h�}����K�j,%  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��0�K�j)%  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���K�h�)��}�(h�Kh�Kh�}����K�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����K�jV%  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjS%  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����K�jS%  sh�Kh�h�h�h�)��}�(h�}��P�K�jt%  sh�K h�h�j  Njd  h�)��}�(h�}�� �K�jw%  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��P�K�jt%  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�@�K�h�)��}�(h�Kh�Kh�}����K�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����K�j�%  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�%  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��@�K�j�%  sh�Kh�h�h�h�)��}�(h�}���K�j�%  sh�K h�h�j  Njd  h�)��}�(h�}��P�K�j�%  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���K�j�%  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���K�h�)��}�(h�Kh�Kh�}�� �K�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� �K�j�%  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�%  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����K�j�%  sh�Kh�h�h�h�)��}�(h�}���K�j
&  sh�K h�h�j  Njd  h�)��}�(h�}�� �K�j&  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���K�j
&  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�p�K�h�)��}�(h�Kh�Kh�}��P�9�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��P�9�j7&  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj4&  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��p�K�j4&  sh�Kh�h�h�h�)��}�(h�}����K�jU&  sh�K h�h�j  Njd  h�)��}�(h�}����K�jX&  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}����K�jU&  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���N�h�)��}�(h�Kh�Kh�}���N�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���N�j�&  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj&  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����N�j&  sh�Kh�h�h�h�)��}�(h�}��ЬN�j�&  sh�K h�h�j  Njd  h�)��}�(h�}����9�j�&  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��ЬN�j�&  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���N�h�)��}�(h�Kh�Kh�}���N�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���N�j�&  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�&  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����N�j�&  sh�Kh�h�h�h�)��}�(h�}��P�N�j�&  sh�K h�h�j  Njd  h�)��}�(h�}��ЩN�j�&  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��P�N�j�&  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� �N�h�)��}�(h�Kh�Kh�}����N�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����N�j'  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj'  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� �N�j'  sh�Kh�h�h�h�)��}�(h�}��P�N�j6'  sh�K h�h�j  Njd  h�)��}�(h�}��`�N�j9'  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��P�N�j6'  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�0�N�h�)��}�(h�Kh�Kh�}����N�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����N�jc'  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj`'  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��0�N�j`'  sh�Kh�h�h�h�)��}�(h�}���N�j�'  sh�K h�h�j  Njd  h�)��}�(h�}����N�j�'  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���N�j�'  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���N�h�)��}�(h�Kh�Kh�}��0�N�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��0�N�j�'  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�'  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����N�j�'  sh�Kh�h�h�h�)��}�(h�}��`�N�j�'  sh�K h�h�j  Njd  h�)��}�(h�}��P�N�j�'  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��`�N�j�'  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� �N�h�)��}�(h�Kh�Kh�}�� �N�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}�� �N�j�'  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�'  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� �N�j�'  sh�Kh�h�h�h�)��}�(h�}����N�j(  sh�K h�h�j  Njd  h�)��}�(h�}��@�N�j(  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}����N�j(  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�O�h�)��}�(h�Kh�Kh�}���O�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���O�jD(  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjA(  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��O�jA(  sh�Kh�h�h�h�)��}�(h�}��PO�jb(  sh�K h�h�j  Njd  h�)��}�(h�}����N�je(  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��PO�jb(  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��O�h�)��}�(h�Kh�Kh�}��`O�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��`O�j�(  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�(  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���O�j�(  sh�Kh�h�h�h�)��}�(h�}���O�j�(  sh�K h�h�j  Njd  h�)��}�(h�}���O�j�(  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���O�j�(  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��O�h�)��}�(h�Kh�Kh�}���O�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���O�j�(  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�(  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���O�j�(  sh�Kh�h�h�h�)��}�(h�}��0O�j�(  sh�K h�h�j  Njd  h�)��}�(h�}��@O�j�(  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��0O�j�(  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��O�h�)��}�(h�Kh�Kh�}���O�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���O�j%)  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj")  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���O�j")  sh�Kh�h�h�h�)��}�(h�}��pO�jC)  sh�K h�h�j  Njd  h�)��}�(h�}��pO�jF)  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��pO�jC)  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��O�h�)��}�(h�Kh�Kh�}���O�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���O�jp)  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjm)  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���O�jm)  sh�Kh�h�h�h�)��}�(h�}���O�j�)  sh�K h�h�j  Njd  h�)��}�(h�}���O�j�)  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���O�j�)  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub��O�h�)��}�(h�Kh�Kh�}���O�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���O�j�)  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�)  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}���O�j�)  sh�Kh�h�h�h�)��}�(h�}��@O�j�)  sh�K h�h�j  Njd  h�)��}�(h�}�� O�j�)  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��@O�j�)  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub�pO�h�)��}�(h�Kh�Kh�}���O�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}���O�j*  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj*  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}��pO�j*  sh�Kh�h�h�h�)��}�(h�}��O�j$*  sh�K h�h�j  Njd  h�)��}�(h�}���O�j'*  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��O�j$*  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub� O�h�)��}�(h�Kh�Kh�}��pN�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}��pN�jQ*  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyjN*  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}�� O�jN*  sh�Kh�h�h�h�)��}�(h�}���O�jo*  sh�K h�h�j  Njd  h�)��}�(h�}���O�jr*  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���O�jo*  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ub���M�h�)��}�(h�Kh�Kh�}����M�h�)��}�(h�}�h�Kh�h�j�  h�)��}�(h�}����M�j�*  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubhyj�*  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�Kh�h�h�h�)��}�(h�Kh�Kh�}����M�j�*  sh�Kh�h�h�h�)��}�(h�}��`�M�j�*  sh�K h�h�j  Njd  h�)��}�(h�}����M�j�*  sh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��`�M�j�*  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bububj   h�ubuh�Kh�h�j  Njd  h�j+  h%h(K ��h*��R�(KKK��hR�CH������Q@            '�@        ��(\�bt@������B@                      �?�t�bubsh�Kh�h�j�  h�hyj  j�  h%h(K ��h*��R�(KKK��hR�C     '�@������B@     g�@�(\�µv@�t�bubsh�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C �������?      �?�������?)\���(�?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C       �?      �?�������?)\���(�?�t�bub�_originalPosition�h�)��}�(h�}�h�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C       �?      �?�������?)\���(�?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C       �?      �?�������?)\���(�?�t�bub�_aspect�h�_adjustable��box��_anchor��C��_stale_viewlim_x���_stale_viewlim_y���_sharex�N�_sharey�hn�bbox�h�dataLim�h�)��}�(h�}�h�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C         033333ӿ      ~@433333�?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �?��G�zd<�t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C       �      �      ��      ���t�bub�_viewLim�j<	  �
transScale�j$	  �	transAxes�h�transLimits�j*	  �	transData�h�_xaxis_transform�h��_yaxis_transform�jO  �_box_aspect�N�_axes_locator��$mpl_toolkits.axes_grid1.axes_divider��AxesLocator���)��}�(�_axes_divider�jA+  �AxesDivider���)��}�(hrhn�_xref��!mpl_toolkits.axes_grid1.axes_size��AxesX���)��}�(hrhnj+  G?�      �_ref_ax�Nub�_yref�jL+  �AxesY���)��}�(hrhnj+  G?�      jQ+  Nub�_fig�hwh�N�_horizontal�]�(jO+  jL+  �Fixed���)��}��
fixed_size�G?�������sbj[+  )��}�j^+  Ksbe�	_vertical�]�jU+  aj+  j+  j+  N�
_xrefindex�K �
_yrefindex�K �_locator�Nub�_nx�K�_ny�K �_nx1�K�_ny1�Kub�
_colorbars�]��spines��matplotlib.spines��Spines���)��}�(�left�jm+  �Spine���)��}�(hp�hqNhrh�hshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h���_hatch_color�(G?陙����G?陙����G?陙����G?�      t��_fill���_original_edgecolor��.8��
_edgecolor�j�+  �_original_facecolor��none��
_facecolor�(G        G        G        G        t��
_us_dashes�K N���
_linewidth�G?�      �
_linestyle��solid��_dashoffset�G        �_dashes�N�_antialiased���_hatch�N�	_capstyle��matplotlib._enums��CapStyle����
projecting���R��
_joinstyle�j�+  �	JoinStyle����miter���R��
spine_type�jr+  �axis��matplotlib.axis��YAxis���)��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~js  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h���_remove_overlapping_locs���isDefault_label���major�j�+  �Ticker���)��}�(je+  �matplotlib.ticker��AutoLocator���)��}�(�_nbins�h�
_symmetric���_prune�N�_min_n_ticks�K�_steps�h%h(K ��h*��R�(KK��hR�C(      �?       @      @      @      $@�t�b�_extended_steps�h%h(K ��h*��R�(KK
��hR�CP�������?�������?      �?      �?      �?       @      @      @      $@      4@�t�b�_integer��j�+  j�+  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~j  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  �j�+  �j�+  j�+  �minor�j�+  )��}�(je+  j�+  �NullLocator���)��}�j�+  j�+  sb�
_formatter�j�+  �NullFormatter���)��}�(j�+  j�+  �locs�]�ububh�h�)��}�(h�h�h�}�(�units finalize�}�K �	functools��partial���h�hn�_unit_change_handler���R���R�(j�+  h���}��event��builtins��object���)��sNt�bs�units�}�Khьmatplotlib.lines��Line2D���)��}�(hp�hqNhrhnhshwhyj�  hz�h{�h|�h}Nh~j�  hNh��h��_line0�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�]�j,  a�remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�]�����h���_dashcapstyle�j�+  �butt���R��_dashjoinstyle�j�+  �round���R��_solidjoinstyle�j,  �_solidcapstyle�j�+  j,  ��R��_linestyles�N�
_drawstyle��default�j�+  G?�      �_dashSeq�N�_dashOffset�G        �_us_dashSeq�N�_us_dashOffset�K j�+  �-��	_invalidx���_color��#111111��_marker��matplotlib.markers��MarkerStyle���)��}�(�_marker_function�h�j1,  �_set_nothing���R��
_fillstyle��full�j-,  �None�j`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�C �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubhyj�  )��}�(h�}�h�Kh�h�j  Nub�	_alt_path�N�_alt_transform�N�_snap_threshold�Nj�+  j,  j�+  j,  �_filled��ub�
_markevery�N�_markersize�G@      j�+  ��_markeredgecolor��auto��_markeredgewidth�G        �_markerfacecolor��auto��_markerfacecoloralt�j�+  �	_invalidy���_pickradius�K�
ind_offset�K �_xorig�]�(K Ke�_yorig�]�(K K ej�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C                �t�b�_xy�h%h(K ��h*��R�(KKK��hR�C                       �?        �t�bj`  j8  jr  j5  �	_subslice���	_x_filled�Nub�recache_always���R�suh�h�K��R�h�Nh���(K K�ub�_autolabelpos���label��matplotlib.text��Text���)��}�(hp�hqNhrNhshwhyj%  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  h#�scalar���hRC8333331@���R�j�  G?�      �_text��	Residuals�j+,  �.15��_fontproperties��matplotlib.font_manager��FontProperties���)��}�(�_family�]��
sans-serif�a�_slant��normal��_variant��normal��_weight��normal��_stretch��normal��_size�G@&      �_file�N�_math_fontfamily��
dejavusans�ub�_usetex���_wrap���_verticalalignment��bottom��_horizontalalignment��center��_multialignment�N�	_rotation��vertical��_transform_rotates_text���_bbox_patch�N�	_renderer�N�_linespacing�G?�333333�_rotation_mode��anchor�ub�
offsetText�jw,  )��}�(hp�hqNhrNhshwhyj1  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j�,  hRC�(\���v@���R�j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  �normal�j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  �baseline�j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nub�labelpad�G@      �
pickradius�K�_major_tick_kw�}�(�gridOn���tick1On���tick2On���label1On���label2On��u�_minor_tick_kw�}�(j�,  �j�,  �j�,  �j�,  �j�,  �u�_scale��matplotlib.scale��LinearScale���)���isDefault_majloc���isDefault_majfmt���isDefault_minfmt���isDefault_minloc���	converter�Nj ,  N�label_position�jr+  �offset_text_position�jr+  �zorder�G?�      �
majorTicks�]�(j�+  �YTick���)��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~ji  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h���_loc�j�,  hRC������ٿ���R��_major��j�,  G        �_width�G?�      �	_base_pad�G@      �_labelrotation�j$,  K ���_zorder�G@ z�G��_tickdir��out��_pad�G@      �_tickmarkers�K K���	tick1line�j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  �None�j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j	-  �_set_tickleft���R�j7,  j8,  j-,  K j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C                       �?        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubhyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �       �       �              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j�,  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nub�	tick2line�j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j.-  �_set_tickright���R�j7,  j8,  j-,  Kj`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j�,  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nub�gridline�j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�jK-  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j�,  ��jQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nub�label1�jw,  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j�,  j�,  �−0.4�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  �center_baseline�j�,  �right�j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nub�label2�jw,  )��}�(hp�hqNhrNhshwhyj   hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j�,  j�,  jw-  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC������ɿ���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�-  j-  ��R�j7,  j8,  j-,  K j`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �       �       �              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j�-  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C        �t�bj�  h%h(K ��h*��R�(KK��hR�C������ɿ�t�bjd,  h%h(K ��h*��R�(KKK��hR�C        ������ɿ�t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C        ������ɿ�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�-  j0-  ��R�j7,  j8,  j-,  Kj`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j�-  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}G?�      h~j2  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�j�-  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j�-  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C������ɿ������ɿ�t�bjd,  h%h(K ��h*��R�(KKK��hR�C         ������ɿ      �?������ɿ�t�bj`  jG  jr  jD  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j�-  j�,  �−0.2�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j�-  j�,  j.  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC        ���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j-  j7,  j8,  j-,  K j`  j-  hyj-  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j>.  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C        �t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C                �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C                �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j2-  j7,  j8,  j-,  Kj`  j-  hyj3-  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j>.  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  jN-  j7,  j8,  j-,  h�j`  j:,  hyjO-  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j>.  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C                �t�bjd,  h%h(K ��h*��R�(KKK��hR�C                       �?        �t�bj`  jV  jr  jS  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j>.  j�,  �0.0�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyj   hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j>.  j�,  j�.  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC�������?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j-  j7,  j8,  j-,  K j`  j-  hyj-  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j�.  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C        �t�bj�  h%h(K ��h*��R�(KK��hR�C�������?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C        �������?�t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C        �������?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j2-  j7,  j8,  j-,  Kj`  j-  hyj3-  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j�.  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  jN-  j7,  j8,  j-,  h�j`  j:,  hyjO-  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j�.  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C�������?�������?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C         �������?      �?�������?�t�b�      j`  je  jr  jb  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j�.  j�,  �0.2�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyj   hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j�.  j�,  j3/  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC�������?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j-  j7,  j8,  j-,  K j`  j-  hyj-  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  jR/  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C        �t�bj�  h%h(K ��h*��R�(KK��hR�C�������?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C        �������?�t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C        �������?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j2-  j7,  j8,  j-,  Kj`  j-  hyj3-  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  jR/  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  jN-  j7,  j8,  j-,  h�j`  j:,  hyjO-  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  jR/  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C�������?�������?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C         �������?      �?�������?�t�bj`  jt  jr  jq  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  jR/  j�,  �0.4�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyj   hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  jR/  j�,  j�/  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC333333�?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j-  j7,  j8,  j-,  K j`  j-  hyj-  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j�/  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C        �t�bj�  h%h(K ��h*��R�(KK��hR�C333333�?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C        333333�?�t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C        333333�?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j2-  j7,  j8,  j-,  Kj`  j-  hyj3-  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j�/  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  jN-  j7,  j8,  j-,  h�j`  j:,  hyjO-  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j�/  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C333333�?333333�?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C         333333�?      �?333333�?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j�/  j�,  �0.6�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyj   hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j�/  j�,  jG0  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC�������?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j-  j7,  j8,  j-,  K j`  j-  hyj-  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  jf0  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j2-  j7,  j8,  j-,  Kj`  j-  hyj3-  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  jf0  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  jN-  j7,  j8,  j-,  h�j`  j:,  hyjO-  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  jf0  ��jQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  jf0  j�,  �0.8�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyj   hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  jf0  j�,  j�0  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubube�
minorTicks�]�j�,  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~j}  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  K j�,  �j�,  G        j�,  G?�      j�,  G@333333j�,  j$,  K ��j�,  Kj�,  j�,  j�,  G@333333j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�0  j-  ��R�j7,  j8,  j-,  K j`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �       �       �              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  KjR,  KjS,  K jT,  ]�K ajV,  ]�K ajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j1  j0-  ��R�j7,  j8,  j-,  Kj`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  KjR,  KjS,  K jT,  ]�KajV,  ]�K ajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�j1  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  ]�(K K ejQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj'  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  K j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyj.  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  K j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububaububj�+  j�+  �ScalarFormatter���)��}�(�_offset_threshold�K�offset�K �
_useOffset��j�,  ��_useMathText���orderOfMagnitude�K �format��%1.1f��_scientific���_powerlimits�]�(J����Ke�
_useLocale��j�+  j�+  j�+  h%h(K ��h*��R�(KK��hR�C8������ٿ������ɿ        �������?�������?333333�?�������?�t�bububj�+  j�+  h�h�)��}�(h�h�h�}�(j�+  }�K j�+  h�h�j�+  ��R���R�(js1  h���}�j�+  j�+  )��sNt�bsj ,  }�Kh�j,  )��}�(hp�hqNhrh�hshwhyjO  hz�h{�h|�h}Nh~j�*  hNh��h��_line0�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�]�j{1  a�remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j,,  j-,  j0,  )��}�(j3,  h�j�1  j4,  ��R�j7,  j8,  j-,  j9,  j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jQ,  �jR,  KjS,  K jT,  ]�(K KejV,  ]�(K K ej�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C                �t�bjd,  h%h(K ��h*��R�(KKK��hR�C                       �?        �t�bj`  j�  jr  j�  jk,  �jl,  Nubjm,  ��R�suh�h�K��R�h�Nh���(K K�ubjs,  �jt,  jw,  )��}�(hp�hqNhrNhshwhyj�	  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�,  hRC    �@���R�j�  G?�      j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@&      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  j�,  j�,  �j�,  Nj�,  Nj�,  G?�333333j�,  j�,  ubj�,  jw,  )��}�(hp�hqNhrNhshwhyj�	  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j�,  hRC�(\���v@���R�j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj�,  G@      j�,  Kj�,  }�(j�,  �j�,  �j�,  �j�,  �j�,  �uj�,  }�(j�,  �j�,  �j�,  �j�,  �j�,  �uj�,  j�,  j�,  �j�,  �j�,  �j�,  �j�,  Nj ,  Nj�,  jr+  j�,  jr+  j�,  G?�      j�,  ]�(j�,  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC������ٿ���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�1  j-  ��R�j7,  j8,  j-,  K j`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �       �       �              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j�1  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j	2  j0-  ��R�j7,  j8,  j-,  Kj`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j�1  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�j$2  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j�1  ��jQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj_  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j�1  j�,  �−0.4�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjf  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j�1  j�,  jO2  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~jH  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC������ɿ���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j}2  j-  ��R�j7,  j8,  j-,  K j`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �       �       �              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  jn2  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�2  j0-  ��R�j7,  j8,  j-,  Kj`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  jn2  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C������ɿ�t�bjd,  h%h(K ��h*��R�(KKK��hR�C      �?������ɿ�t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C      �?������ɿ�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�j�2  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  jn2  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C������ɿ������ɿ�t�bjd,  h%h(K ��h*��R�(KKK��hR�C         ������ɿ      �?������ɿ�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyjL  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  jn2  j�,  �−0.2�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjR  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  jn2  j�,  j�2  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC        ���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�1  j7,  j8,  j-,  K j`  j-  hyj�1  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j3  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j2  j7,  j8,  j-,  Kj`  j-  hyj2  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j3  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C      �?        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C      �?        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j'2  j7,  j8,  j-,  h�j`  j:,  hyj(2  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j3  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C                �t�bjd,  h%h(K ��h*��R�(KKK��hR�C                       �?        �t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj_  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j3  j�,  �0.0�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjf  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j3  j�,  j~3  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC�������?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�1  j7,  j8,  j-,  K j`  j-  hyj�1  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j�3  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j2  j7,  j8,  j-,  Kj`  j-  hyj2  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j�3  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C�������?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C      �?�������?�t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C      �?�������?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j'2  j7,  j8,  j-,  h�j`  j:,  hyj(2  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j�3  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C�������?�������?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C         �������?      �?�������?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj_  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j�3  j�,  �0.2�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjf  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j�3  j�,  j4  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC�������?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�1  j7,  j8,  j-,  K j`  j-  hyj�1  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j'4  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j2  j7,  j8,  j-,  Kj`  j-  hyj2  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j'4  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C�������?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C      �?�������?�t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C      �?�������?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j'2  j7,  j8,  j-,  h�j`  j:,  hyj(2  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j'4  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C�������?�������?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C         �������?      �?�������?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj_  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j'4  j�,  �0.4�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjf  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j'4  j�,  j�4  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC333333�?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�1  j7,  j8,  j-,  K j`  j-  hyj�1  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j�4  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j2  j7,  j8,  j-,  Kj`  j-  hyj2  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j�4  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C333333�?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C      �?333333�?�t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C      �?333333�?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j'2  j7,  j8,  j-,  h�j`  j:,  hyj(2  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j�4  ��jQ,  �j�  h%h(K ��h*��R�(KK��hR�C              �?�t�bj�  h%h(K ��h*��R�(KK��hR�C333333�?333333�?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C         333333�?      �?333333�?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj_  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j�4  j�,  �0.6�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjf  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j�4  j�,  j5  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�,  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC�������?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�1  j7,  j8,  j-,  K j`  j-  hyj�1  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�K ajV,  j;5  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j2  j7,  j8,  j-,  Kj`  j-  hyj2  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  ]�KajV,  j;5  ��jQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j'2  j7,  j8,  j-,  h�j`  j:,  hyj(2  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  j;5  ��jQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj_  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  j;5  j�,  �0.8�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjf  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j;5  j�,  j�5  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububej�0  ]�j�,  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  K j�,  �j�,  G        j�,  G?�      j�,  G@333333j�,  j$,  K ��j�,  Kj�,  j�,  j�,  G@333333j�,  K K��j�,  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�5  j-  ��R�j7,  j8,  j-,  K j`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �       �       �              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  KjR,  KjS,  K jT,  ]�K ajV,  ]�K ajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�5  j0-  ��R�j7,  j8,  j-,  Kj`  j-  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  KjR,  KjS,  K jT,  ]�KajV,  ]�K ajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyjO  hz�h{�h|�h}G?�      h~j  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�j�5  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K KejV,  ]�(K K ejQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyjs  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  K j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjz  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  K j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  jz-  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububaubj�,  G@      �_bounds�Nhٌoutward�G        ��j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C         �G�zֿ        �p=
ף�?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ub�_patch_type��line��_patch_transform�j�  )��}�(h�}�h�Kh�h�j  Nububj{-  jt+  )��}�(hp�hqNhrh�hshwhyjO  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  j�+  j�+  �j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  K N��j�+  G?�      j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j�+  j�+  j�+  j�+  j{-  j�+  j�+  j�,  G@      j-6  Nh�j/6  j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C       �?�G�zֿ      �?�p=
ף�?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubj86  j96  j:6  j�  )��}�(h�}�h�Kh�h�j  Nububj�,  jt+  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  j�+  j�+  �j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  K N��j�+  G?�      j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j�+  j�+  j�+  j�+  j�,  j�+  j�+  �XAxis���)��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~j�	  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  �j�+  �j�+  j�+  )��}�(je+  j�+  )��}�(j�+  hj�+  �j�+  Nj�+  Kj�+  h%h(K ��h*��R�(KK��hR�C(      �?       @      @      @      $@�t�bj�+  h%h(K ��h*��R�(KK
��hR�CP�������?�������?      �?      �?      �?       @      @      @      $@      4@�t�bj�+  �j�+  je6  ubj�+  jZ1  )��}�(j]1  Kj^1  K j_1  �j�,  �j`1  �ja1  K jb1  �%1.0f�jd1  �je1  jf1  jg1  �j�+  je6  j�+  h%h(K ��h*��R�(KK��hR�C             @@     @�@�t�bububj�+  j�+  )��}�(je+  j�+  )��}�j�+  je6  sbj�+  j�+  )��}�(j�+  je6  j�+  ]�ububh�h�)��}�(h�h�h�}�(j�+  }�K j�+  h�h�j�+  ��R���R�(j�6  h���}�j�+  j�+  )��sNt�bsj ,  }�Kh�j{1  jm,  ��R�suh�h�K��R�h�Nh���(K K�ubjs,  �jt,  jw,  )��}�(hp�hqNhrNhshwhyj{	  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  G?�      j�  j�,  hRC4333331@���R�j�,  �Distribution�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@&      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  �top�j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj�,  jw,  )��}�(hp�hqNhrNhshwhyj�	  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j�,  hRC4333332@���R�j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj�,  G@      j�,  Kj�,  }�(j�,  �j�,  �j�,  �j�,  �j�,  �uj�,  }�(j�,  �j�,  �j�,  �j�,  �j�,  �uj�,  j�,  )��j�,  �j�,  �j�,  �j�,  �j�,  Nj ,  Nj�,  j�,  j�,  j�,  j�,  G?�      j�,  ]�(j�+  �XTick���)��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~j�	  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC        ���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�6  �_set_tickdown���R�j7,  j8,  j-,  Kj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C        �               �      �?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubhyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                       �      �       �                      �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�6  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�C        �t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C                �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C                �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j(7  �_set_tickup���R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�6  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}G?�      h~j8
  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�jD7  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j�6  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj8  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�6  j�  K j�,  �0�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjE  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�6  j�  Kj�,  jo7  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~jw
  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC     @@���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�7  j�6  ��R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                       �      �       �                      �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�7  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�C     @@�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C     @@        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C     @@        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�7  j*7  ��R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�7  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}G?�      h~j�
  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�j�7  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j�7  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�7  j�  K j�,  �500�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyj1  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�7  j�  Kj�,  j8  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC     @�@���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�6  j7,  j8,  j-,  Kj`  j�6  hyj�6  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j78  ��jV,  ]�K ajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j,7  j7,  j8,  j-,  Kj`  j�6  hyj-7  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j78  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}G?�      h~j8
  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  jG7  j7,  j8,  j-,  h�j`  j:,  hyjH7  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j78  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj8  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j78  j�  K j�,  �1000�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjE  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j78  j�  Kj�,  j�8  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububej�0  ]�j�6  )��}�(hp�hqNhrh�hshwhyNhz�h{�h|�h}Nh~j�
  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  K j�,  �j�,  G        j�,  G?�      j�,  G@333333j�,  j$,  K ��j�,  Kj�,  j�,  j�,  G@333333j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�8  j�6  ��R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                       �      �       �                      �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  KjR,  KjS,  K jT,  ]�K ajV,  ]�K ajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�8  j*7  ��R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  KjR,  KjS,  K jT,  ]�K ajV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}G?�      h~j4  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�j�8  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K K ejV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  K j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyj	  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  Kj�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububa�_tick_position�j�,  ubj�,  G@      j-6  Nh�j/6  j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C                      �@        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubj86  j96  j:6  j�  )��}�(h�}�h�Kh�h�j  Nububj�6  jt+  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  j�+  j�+  �j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  K N��j�+  G?�      j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j�+  j�+  j�+  j�+  j�6  j�+  je6  j�,  G@      j-6  Nh�j/6  j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C               �?     �@      �?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubj86  j96  j:6  j�  )��}�(h�}�h�Kh�h�j  Nububub�xaxis�je6  �yaxis�j�+  j�+  �white��_frameon���
_axisbelow���_rasterization_zorder�N�ignore_existing_data_limits��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ub�_autoscaleXon���_autoscaleYon���_xmargin�G?��������_ymargin�G?��������_tight�N�_use_sticky_edges���
_get_lines��matplotlib.axes._base��_process_plot_var_args���)��}�(�axes�hǌcommand��plot�ub�_get_patches_for_fill�jc9  )��}�(jf9  h�jg9  �fill�ub�_gridOn���lines�j�1  �patches�]�(�matplotlib.patches��	Rectangle���)��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jP  hNh��h��
_nolegend_�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  (G        G        G        G?�      t�j�+  �j�+  Nj�+  j�+  j�+  h%h(K ��h*��R�(KK��hR�C �?�������?TTTTTT�?      �?�t�bj�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  �_x0�j�9  �_y0�j�,  hRC      �����R�j�,  j�,  hRC      @���R��_height�j�,  hRC��G�zd<���R��angle�G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�9  j�9  j�,  hRC���Q������R�j�,  j�,  hRC        ���R�j�9  j�,  hRCp�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�9  j�9  j�,  hRCq=
ףp�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j1  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�9  j�9  j�,  hRC)\���(�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j|  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j:  j�9  j�,  hRC�z�G᪼���R�j�,  j�,  hRC        ���R�j�9  j�,  hRCp�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j:  j�9  j�,  hRC�����������R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j<:  j�9  j�,  hRCR���Q�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j]  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jY:  j�9  j�,  hRC
ףp=
�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jv:  j�9  j�,  hRC��(\�¥����R�j�,  j�,  hRC        ���R�j�9  j�,  hRCp�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�:  j�9  j�,  hRC{�G�z�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j>  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�:  j�9  j�,  hRC433333�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRCp�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�:  j�9  j�,  hRC�Q��롼���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�:  j�9  j�,  hRC�p=
ף�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j;  j�9  j�,  hRC���Q������R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jj  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j$;  j�9  j�,  hRC(\���(�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRCp�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jA;  j�9  j�,  hRC�����������R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j   hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j^;  j�9  j�,  hRC
ףp=
�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jK  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j{;  �      j�9  j�,  hRCz�G�z�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRCp�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�;  j�9  j�,  hRC�Q��둼���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�;  j�9  j�,  hRC���Q������R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j,  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�;  j�9  j�,  hRC�����������R�j�,  j�,  hRC        ���R�j�9  j�,  hRCp�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jw  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�;  j�9  j�,  hRC|�G�z�����R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j<  j�9  j�,  hRC���Q�~����R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j)<  j�9  j�,  hRCx�G�zt����R�j�,  j�,  hRC        ���R�j�9  j�,  hRCp�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jX  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jF<  j�9  j�,  hRC��G�zd����R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jc<  j�9  j�,  hRC        ���R�j�,  j�,  hRC      ~@���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�<  j�9  j�,  hRC��G�zd<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j9  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�<  j�9  j�,  hRC��G�zt<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�<  j�9  j�,  hRC���Q�~<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC`�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�<  j�9  j�,  hRCx�G�z�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�<  j�9  j�,  hRC�������<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~je  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j=  j�9  j�,  hRC���Q��<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j.=  j�9  j�,  hRC�Q���<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jK=  j�9  j�,  hRC|�G�z�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jF  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jh=  j�9  j�,  hRCףp=
�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�=  j�9  j�,  hRC�������<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC`�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�=  j�9  j�,  hRC(\���(�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j'  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�=  j�9  j�,  hRC���Q��<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jr  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�=  j�9  j�,  hRC�p=
ף�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�=  j�9  j�,  hRC�Q���<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j>  j�9  j�,  hRC433333�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jS  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j3>  j�9  j�,  hRC|�G�z�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC`�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jP>  j�9  j�,  hRC��(\�¥<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jm>  j�9  j�,  hRC
ףp=
�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j4  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�>  j�9  j�,  hRCR���Q�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�>  j�9  j�,  hRC�������<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�>  j�9  j�,  hRC�z�G�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�>  j�9  j�,  hRC*\���(�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC`�G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j`  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�>  j�9  j�,  hRCp=
ףp�<���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j�9  j�+  (G?�G?ܜ�����G?�TTTTTTG?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j?  j�9  j�,  hRC���Q��<���R�j�,  j�,  hRC     �L@���R�j�9  j�,  hRC��G�zd<���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  h%h(K ��h*��R�(KK��hR�C �������?xxxxxx�?�������?      �?�t�bj�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j8?  j�9  j�,  hRC033333ӿ���R�j�,  j�,  hRC      �?���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jA  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j[?  j�9  j�,  hRC<5^�Iҿ���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC0�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jx?  j�9  j�,  hRCI7�A`�п���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�?  j�9  j�,  hRC�rh��|Ͽ���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j"  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�?  j�9  j�,  hRC�v��/Ϳ���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jm  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�?  j�9  j�,  hRC�z�G�ʿ���R�j�,  j�,  hRC       @���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�?  j�9  j�,  hRC�~j�t�ȿ���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j	@  j�9  j�,  hRC��ʡEƿ���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jN  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j&@  j�9  j�,  hRC&����ÿ���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jC@  j�9  j�,  hRC>�l��������R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j`@  j�9  j�,  hRC���Q������R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j/  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j}@  j�9  j�,  hRC�&1������R�j�,  j�,  hRC      5@���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jz  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�@  j�9  j�,  hRC/�$������R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�@  j�9  j�,  hRC@7�A`尿���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j   hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�@  j�9  j�,  hRC�~j�t������R�j�,  j�,  hRC        ���R�j�9  j�,  hRC0�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j[   hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�@  j�9  j�,  hRC���Q������R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�   hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jA  j�9  j�,  hRC�~j�t������R�j�,  j�,  hRC     �P@���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�   hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j+A  j�9  j�,  hRC�j�t�x?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC0�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j<!  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jHA  j�9  j�,  hRC j�t��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�!  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jeA  j�9  j�,  hRC0/�$��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�!  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�A  j�9  j�,  hRC���Q��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC0�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j"  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�A  j�9  j�,  hRC4�����?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jh"  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�A  j�9  j�,  hRCj�t��?���R�j�,  j�,  hRC      4@���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�"  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�A  j�9  j�,  hRC�v��/�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC0�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�"  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�A  j�9  j�,  hRCP7�A`��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jI#  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jB  j�9  j�,  hRC833333�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�#  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j0B  j�9  j�,  hRC /�$��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�#  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jMB  j�9  j�,  hRC+����?���R�j�,  j�,  hRC      0@���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j*$  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jjB  j�9  j�,  hRC�&1��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC �O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~ju$  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�B  j�9  j�,  hRC�"��~j�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�$  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�B  j�9  j�,  hRC���Q��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j%  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�B  j�9  j�,  hRCR��n��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jV%  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�B  j�9  j�,  hRCF�l����?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�%  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�B  j�9  j�,  hRC:�A`���?���R�j�,  j�,  hRC      @���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�%  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jC  j�9  j�,  hRC.�����?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j7&  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j5C  j�9  j�,  hRC"��Q��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC �O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�&  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jRC  j�9  j�,  hRC��ʡE�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�&  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  joC  j�9  j�,  hRC��C�l�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j'  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�C  j�9  j�,  hRC�~j�t��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jc'  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�C  j�9  j�,  hRC�|?5^��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�'  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�C  j�9  j�,  hRC�z�G��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�'  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�C  j�9  j�,  hRC�x�&1�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC �O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jD(  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j D  j�9  j�,  hRC�v��/�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�(  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jD  j�9  j�,  hRC�t�V�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�(  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j:D  j�9  j�,  hRC�rh��|�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j%)  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jWD  j�9  j�,  hRCS���Q�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jp)  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  jtD  j�9  j�,  hRCM7�A`��?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j�)  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�D  j�9  j�,  hRCH����x�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC �O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~j*  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�D  j�9  j�,  hRC@5^�I�?���R�j�,  j�,  hRC        ���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ubjs9  )��}�(hp�hqNhrh�hshwhyh�hz�h{�h|�h}Nh~jQ*  hNh��h�jv9  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jp9  �remove���R�h�Nh�Nh�Nh�Nh�h�h�h�]�j�,  hRC        ���R�a]�����h��j�+  j�9  j�+  �j�+  Nj�+  j�+  j�+  j>?  j�+  (G?�������G?�xxxxxxG?�������G?�      t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  j�D  j�9  j�,  hRC:��v���?���R�j�,  j�,  hRC      �?���R�j�9  j�,  hRC@�O��n�?���R�j�9  G        ube�texts�]��tables�]��artists�]��images�]��_mouseover_set�h��_OrderedSet���)��}��_od��collections��OrderedDict���)R�sb�
child_axes�]��_current_image�N�_projection_init�N�legend_�Nj�D  ]��
containers�]�(�matplotlib.container��BarContainer���(jt9  j�9  j�9  j�9  j�9  j:  j.:  jK:  jh:  j�:  j�:  j�:  j�:  j�:  j;  j3;  jP;  jm;  j�;  j�;  j�;  j�;  j�;  j<  j8<  jU<  jr<  j�<  j�<  j�<  j�<  j=  j =  j==  jZ=  jw=  j�=  j�=  j�=  j�=  j>  j%>  jB>  j_>  j|>  j�>  j�>  j�>  j�>  j?  t�����}�(jo9  ]�(jt9  j�9  j�9  j�9  j�9  j:  j.:  jK:  jh:  j�:  j�:  j�:  j�:  j�:  j;  j3;  jP;  jm;  j�;  j�;  j�;  j�;  j�;  j<  j8<  jU<  jr<  j�<  j�<  j�<  j�<  j=  j =  j==  jZ=  jw=  j�=  j�=  j�=  j�=  j>  j%>  jB>  j_>  j|>  j�>  j�>  j�>  j�>  j?  e�errorbar�N�
datavalues�h%h(K ��h*��R�(KK2��hR�B�        @                                                                                                                                                                                                      ~@                                                                                                                                                                                             �L@�t�b�orientation��
horizontal�h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�j�D  �remove���R�h��_container0��stale��ubj�D  (j*?  jM?  jj?  j�?  j�?  j�?  j�?  j�?  j@  j5@  jR@  jo@  j�@  j�@  j�@  j�@  j A  jA  j:A  jWA  jtA  j�A  j�A  j�A  j�A  jB  j"B  j?B  j\B  jyB  j�B  j�B  j�B  j�B  j
C  j'C  jDC  jaC  j~C  j�C  j�C  j�C  j�C  jD  j,D  jID  jfD  j�D  j�D  j�D  t�����}�(jo9  ]�(j*?  jM?  jj?  j�?  j�?  j�?  j�?  j�?  j@  j5@  jR@  jo@  j�@  j�@  j�@  j�@  j A  jA  j:A  jWA  jtA  j�A  j�A  j�A  j�A  jB  j"B  j?B  j\B  jyB  j�B  j�B  j�B  j�B  j
C  j'C  jDC  jaC  j~C  j�C  j�C  j�C  j�C  jD  j,D  jID  jfD  j�D  j�D  j�D  ej�D  Nj�D  h%h(K ��h*��R�(KK2��hR�B�        �?                                       @                                              5@                                     �P@                                              4@                                      0@                                              @                                                                                                                              �?�t�bjE  jE  h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�j�D  �remove���R�h��_container1�jE  �ube�_autotitlepos���title�jw,  )��}�(hp�hqNhrh�hshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  G?�      j�  G?�      j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  �normal�j�,  j�,  j�,  G@(      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nub�_left_title�jw,  )��}�(hp�hqNhrh�hshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  G        j�  G?�      j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j6E  j�,  j�,  j�,  G@(      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nub�_right_title�jw,  )��}�(hp�hqNhrh�hshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  G?�      j�  G?�      j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j6E  j�,  j�,  j�,  G@(      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nub�titleOffsetTrans�j�  �patch�js9  )��}�(hp�hqNhrNhshwhyh�hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  j�+  j�+  �j�+  j-  j�+  j�+  j�+  jO9  j�+  (G?�      G?�      G?�      G?�      t�j�+  K N��j�+  G        j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  G        j�9  G        j�,  G?�      j�9  G?�      j�9  G        ub�axison���	fmt_xdata�N�	fmt_ydata�N�	_navigate���_navigate_mode�N�_shared_x_axes�N�_shared_y_axes�]�(h�hne�_twinned_axes�Nub��e�_default�N�_ind�Kubj�D  ]�jn9  ]�jo9  ]�j�D  ]�j�D  ]��legends�]��subfigs�]��suppressComposite�Nh�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ub�_canvas_callbacks�h�)��}�(h�h�h�}�(�button_press_event�}��scroll_event�}��key_press_event�}�uh�h�K��R�h�Nh���ub�_button_pick_id�K �_scroll_pick_id�K�bbox_inches�j  �dpi_scale_trans�j  �_dpi�G@R      j!+  j  �figbbox�j  �transFigure�j  �transSubfigure�j  jVE  js9  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  (G?�      G?�      G?�      G        t�j�+  �j�+  j�E  j�+  j�E  j�+  jcE  j�+  (G?�      G?�      G?�      G?�      t�j�+  K N��j�+  G        j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  K j�9  K j�,  Kj�9  Kj�9  G        ub�subplotpars�ht�SubplotParams���)��}�(�validate��jr+  G?�      j�,  G?�      j{-  G?�������j�6  G?�(�\)�wspace�G?ə������hspace�G?ə�����ub�_constrained��j^9  ��_tight_parameters�}��_axstack�h�)��}�(h�Kh�]�(Khǆ�Khn��ejoE  NjpE  Kub�_axobservers�h�)��}�(h�h�h�}��_axes_change_event�}�sh�h�K��R�h�Nh���ub�_cachedRenderer�N�_constrained_layout_pads�}�(�w_pad�G?�U�.r��h_pad�G?�U�.r�j�E  G?�z�G�{j�E  G?�z�G�{u�number�K�__mpl_version__��3.4.3�ubhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�hwh҆�R�h�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��h�j�  j+  h�)��}�(h�}�h�K h�h�j�  h%h(K ��h*��R�(KKK��hR�C       �?      �?�������?)\���(�?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �      ��t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C                       �?      �?�t�bubj+  hj+  j+  j+  j+  j+  �j+  �j+  Nj +  Nj!+  j  j"+  h�)��}�(h�}�h�Kh�h�j�  h%h(K ��h*��R�(KKK��hR�C       �?033333ӿ������@433333�?�t�bj�  h%h(K ��h*��R�(KK��hR�C      �?      �<�t�bj�  �j�  h%h(K ��h*��R�(KKK��hR�C       �      �      ��      ���t�bubj8+  j�  j9+  j�  j:+  j  j;+  j�  j<+  j  j=+  j!  j>+  j�  j?+  Nj@+  jC+  )��}�(jF+  jI+  jf+  K jg+  K jh+  Kji+  Kubjj+  ]�jl+  jo+  )��}�(jr+  jt+  )��}�(hp�hqNhrhnhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  j�+  j�+  �j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  K N��j�+  G?�      j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j�+  j�+  j�+  j�+  jr+  j�+  j�+  j�,  G@      j-6  Nh�j/6  j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C         �G�zֿ        �p=
ף�?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubj86  j96  j:6  j�  )��}�(h�}�h�Kh�h�j  Nububj{-  jt+  )��}�(hp�hqNhrhnhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  j�+  j�+  �j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  K N��j�+  G?�      j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j�+  j�+  j�+  j�+  j{-  j�+  j�+  j�,  G@      j-6  Nh�j/6  j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C       �?�G�zֿ      �?�p=
ף�?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubj86  j96  j:6  j�  )��}�(h�}�h�Kh�h�j  Nububj�,  jt+  )��}�(hp�hqNhrhnhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  j�+  j�+  �j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  K N��j�+  G?�      j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j�+  j�+  j�+  j�+  j�,  j�+  jd6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~j@  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  �j�+  �j�+  j�+  )��}�(je+  j�+  )��}�(j�+  hj�+  �j�+  Nj�+  Kj�+  h%h(K ��h*��R�(KK��hR�C(      �?       @      @      @      $@�t�bj�+  h%h(K ��h*��R�(KK
��hR�CP�������?�������?      �?      �?      �?       @      @      @      $@      4@�t�bj�+  �j�+  j?F  ubj�+  jZ1  )��}�(j]1  Kj^1  K j_1  �j�,  �j`1  �ja1  K jb1  �%1.1f�jd1  �je1  jf1  jg1  �j�+  j?F  j�+  h%h(K ��h*��R�(KK��hR�CX�������?      �?433333�?gfffff�?�������?�������?       @������@433333@������@ffffff@�t�bububj�+  j�+  )��}�(je+  j�+  )��}�j�+  j?F  sbj�+  j�+  )��}�(j�+  j?F  j�+  ]�ububh�h�)��}�(h�h�h�}�(j�+  }�K j�+  h�hnj�+  ��R���R�(jpF  h���}�j�+  j�+  )��sNt�bsj ,  }�Kh�j,  jm,  ��R�suh�h�K��R�h�Nh���(K K�ubjs,  �jt,  jw,  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  G?�      j�  j�,  hRC4333331@���R�j�,  �Predicted Value�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@&      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj�,  jw,  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  Kj�  j�,  hRC4333332@���R�j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj�,  G@      j�,  Kj�,  }�(j�,  �j�,  �j�,  �j�,  �j�,  �uj�,  }�(j�,  �j�,  �j�,  �j�,  �j�,  �uj�,  j�,  )��j�,  �j�,  �j�,  �j�,  �j�,  Nj ,  Nj�,  j�,  j�,  j�,  j�,  G?�      j�,  ]�(j�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC�������?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�F  j�6  ��R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                       �      �       �                      �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�F  ��jV,  ]�K ajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�F  j*7  ��R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�F  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�j�F  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j�F  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj9  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�F  j�  K j�,  �0.8�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjF  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�F  j�  Kj�,  j"G  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~j  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC      �?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�jPG  j�6  ��R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                       �      �       �                      �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  jAG  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�C      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C      �?        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C      �?        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�G  j*7  ��R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  jAG  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~jU  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�j�G  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  jAG  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK��hR�C      �?      �?�t�bj�  h%h(K ��h*��R�(KK��hR�C              �?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C       �?              �?      �?�t�bj`  jd  jr  j]  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj$  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  jAG  j�  K j�,  �1.0�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyj2  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  jAG  j�  Kj�,  j�G  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC433333�?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�G  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�C433333�?�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C433333�?        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C433333�?        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�G  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  h�j`  j:,  hyj�F  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j�G  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK��hR�C433333�?433333�?�t�bj�  h%h(K ��h*��R�(KK��hR�C              �?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C 433333�?        433333�?      �?�t�bj`  j{  jr  jx  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj9  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�G  j�  K j�,  �1.2�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjF  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�G  j�  Kj�,  jQH  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRCgfffff�?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  jpH  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�Cgfffff�?�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�Cgfffff�?        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�Cgfffff�?        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  jpH  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  h�j`  j:,  hyj�F  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  jpH  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK��hR�Cgfffff�?gfffff�?�t�bj�  h%h(K ��h*��R�(KK��hR�C              �?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C gfffff�?        gfffff�?      �?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj9  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  jpH  j�  K j�,  �1.4�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjF  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  jpH  j�  Kj�,  j�H  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC�������?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�H  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�C�������?�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C�������?        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C�������?        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�H  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  h�j`  j:,  hyj�F  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j�H  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK��hR�C�������?�������?�t�bj�  h%h(K ��h*��R�(KK��hR�C              �?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C �������?        �������?      �?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj9  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�H  j�  K j�,  �1.6�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjF  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�H  j�  Kj�,  jeI  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC�������?���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�I  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�C�������?�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C�������?        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C�������?        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�I  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  ��      j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  h�j`  j:,  hyj�F  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j�I  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK��hR�C�������?�������?�t�bj�  h%h(K ��h*��R�(KK��hR�C              �?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C �������?        �������?      �?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj9  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�I  j�  K j�,  �1.8�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjF  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�I  j�  Kj�,  j�I  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC       @���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  jJ  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�C       @�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C       @        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C       @        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  jJ  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  h�j`  j:,  hyj�F  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  jJ  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK��hR�C       @       @�t�bj�  h%h(K ��h*��R�(KK��hR�C              �?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C        @               @      �?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj9  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  jJ  j�  K j�,  �2.0�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjF  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  jJ  j�  Kj�,  jyJ  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC������@���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�J  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�C������@�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C������@        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C������@        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�J  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  h�j`  j:,  hyj�F  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j�J  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK��hR�C������@������@�t�bj�  h%h(K ��h*��R�(KK��hR�C              �?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C ������@        ������@      �?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj9  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�J  j�  K j�,  �2.2�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjF  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�J  j�  Kj�,  jK  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC433333@���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j"K  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�C433333@�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C433333@        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C433333@        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j"K  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  h�j`  j:,  hyj�F  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j"K  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK��hR�C433333@433333@�t�bj�  h%h(K ��h*��R�(KK��hR�C              �?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C 433333@        433333@      �?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj9  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j"K  j�  K j�,  �2.4�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjF  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j"K  j�  Kj�,  j�K  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRC������@���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�K  ��jV,  ]�K ajQ,  �j�  h%h(K ��h*��R�(KK��hR�C������@�t�bj�  h%h(K ��h*��R�(KK��hR�C        �t�bjd,  h%h(K ��h*��R�(KKK��hR�C������@        �t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C������@        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j�K  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  h�j`  j:,  hyj�F  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j�K  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK��hR�C������@������@�t�bj�  h%h(K ��h*��R�(KK��hR�C              �?�t�bjd,  h%h(K ��h*��R�(KKK��hR�C ������@        ������@      �?�t�bj`  j�  jr  j�  jk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj9  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�K  j�  K j�,  �2.6�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjF  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j�K  j�  Kj�,  jL  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububj�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  j�,  hRCffffff@���R�j�,  �j�,  G        j�,  G?�      j�,  G@      j�,  j$,  K ��j�,  G@ z�G�j�,  j�,  j�,  G@      j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j6L  ��jV,  ]�K ajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  Kj`  j�6  hyj�F  jE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  G@ z�G�jR,  KjS,  K jT,  j6L  ��jV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  j�F  j7,  j8,  j-,  h�j`  j:,  hyj�F  jE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  j6L  ��jV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyj9  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j6L  j�  K j�,  �2.8�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjF  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  j6L  j�  Kj�,  j�L  j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububej�0  ]�j�6  )��}�(hp�hqNhrhnhshwhyNhz�h{�h|�h}Nh~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�,  K j�,  �j�,  G        j�,  G?�      j�,  G@333333j�,  j$,  K ��j�,  Kj�,  j�,  j�,  G@333333j�,  KK��j�,  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�L  j�6  ��R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                       �      �       �                      �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  KjR,  KjS,  K jT,  ]�K ajV,  ]�K ajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj!-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j-  j*,  �j+,  j�,  j-,  j0,  )��}�(j3,  h�j�L  j*7  ��R�j7,  j8,  j-,  Kj`  j�6  hyj  )��}�(h�}�h�Kh�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubjE,  NjF,  NjG,  G?�      j�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G        j�+  �jK,  j�,  jM,  G?�      jN,  jO,  jP,  j�+  j�,  KjR,  KjS,  K jT,  ]�K ajV,  ]�KajQ,  �j�  Nj�  Njd,  Nj`  Njr  Njk,  �jl,  Nubj>-  j,  )��}�(hp�hqNhrNhshwhyj!  hz�h{�h|�h}G?�      h~j�  hNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j,  j,  j,  j,  j,  j,  j,  j!,  j",  Nj#,  j$,  j�+  G?�      j%,  Nj&,  G        j',  Nj(,  K j�+  j),  j*,  �j+,  j�+  j-,  j0,  )��}�(j3,  h�j�L  j4,  ��R�j7,  j8,  j-,  h�j`  j:,  hyj�  )��}�(h�}�h�Kh�h�j  NubjE,  NjF,  NjG,  Nj�+  j,  j�+  j,  jH,  �ubjI,  NjJ,  G@      j�+  �jK,  jL,  jM,  G        jN,  jO,  jP,  j�+  jR,  KjS,  K jT,  ]�(K K ejV,  ]�(K KejQ,  �j�  h%h(K ��h*��R�(KK ��hR�j@,  t�bj�  h%h(K ��h*��R�(KK ��hR�j@,  t�bjd,  h%h(K ��h*��R�(KK K��hR�j@,  t�bj`  jc  )��}�(jf  h%h(K ��h*��R�(KK K��hR�j@,  t�bjm  Njn  K�jo  G?�q�q��jp  �jq  �ubjr  Njk,  �jl,  Nubjj-  jw,  )��}�(hp�hqNhrNhshwhyjM  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  K j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�6  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj|-  jw,  )��}�(hp�hqNhrNhshwhyjT  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  Kj�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j�,  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nububaj)9  j�,  ubj�,  G@      j-6  Nh�j/6  j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C p=
ףp�?        q=
ףp@        �t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubj86  j96  j:6  j�  )��}�(h�}�h�Kh�h�j  Nububj�6  jt+  )��}�(hp�hqNhrhnhshwhyj!  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  j�+  j�+  �j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  K N��j�+  G?�      j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j�+  j�+  j�+  j�+  j�6  j�+  j?F  j�,  G@      j-6  Nh�j/6  j`  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�C p=
ףp�?      �?q=
ףp@      �?�t�bjm  Njn  Kjo  G?�q�q��jp  �jq  �ubj86  j96  j:6  j�  )��}�(h�}�h�Kh�h�j  NubububjM9  j?F  jN9  j�+  j�+  jO9  jP9  �jQ9  �jR9  NjS9  �h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubjZ9  �j[9  �j\9  G?�������j]9  G?�������j^9  Nj_9  �j`9  jc9  )��}�(jf9  hnjg9  jh9  ubji9  jc9  )��}�(jf9  hnjg9  jl9  ubjm9  �jn9  j,  jo9  ]�j�D  ]�j�D  ]�j�D  ]�j�D  ]�j�D  j�D  )��}�j�D  j�D  )R�sbj�D  ]�j�D  Nj�D  hl}���j�D  �matplotlib.legend��Legend���)��}�(hp�hqNhrhnhshwhyj�  )��}�(h�}�h�Kh�h�j  Nubhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�hn�_remove_legend���R�h�Nh�Nh�Nh�Nh�h�h�h�]�]�����h���prop�j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ub�	_fontsize�G@$      j�D  ]�(jw,  )��}�(hp�hqNhrNhshwhyhڌCompositeAffine2D���)��}�(h�Kh�Kh�}�h�K h�h�j  Nh�j  )��}�(h�}���N�j~M  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?        �p=
�#�@              �?*\���hu@                      �?�t�bubj   j  )��}�(h�}���N�j~M  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?        �p=
�#�@              �?*\���hu@                      �?�t�bubhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  K j�,  �Train $R^2 = 1.000$�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubjw,  )��}�(hp�hqNhrNhshwhyj}M  )��}�(h�Kh�Kh�}�h�K h�h�j  Nh�j  )��}�(h�}��`N�j�M  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?        �p=
�#�@              �?]���(<t@                      �?�t�bubj   j  )��}�(h�}��`N�j�M  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?        �p=
�#�@              �?]���(<t@                      �?�t�bubhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  K j�,  �Test $R^2 = 0.945$�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@$      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nube�legendHandles�]�(js9  )��}�(hp�hqNhrhnhshwhyj}M  )��}�(h�Kh�Kh�}�h�K h�h�j  Nh�j  )��}�(h�}��@N�j�M  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}��@N�j�M  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?        �p=
�C�@              �?*\���hu@                      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?        �p=
�C�@              �?*\���hu@                      �?�t�bubhz�h{�h|�h}Nh~NhNh��h�j�M  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  (G?�G?ܜ�����G?�TTTTTTKt�j�+  �j�+  �b�j�+  j�M  j�+  j�M  j�+  j�M  j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  G�       j�9  G�       j�,  G@4      j�9  G@      j�9  G        ubjs9  )��}�(hp�hqNhrhnhshwhyj}M  )��}�(h�Kh�Kh�}�h�K h�h�j  Nh�j  )��}�(h�}���N�j�M  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}���N�j�M  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?        �p=
�C�@              �?]���(<t@                      �?�t�bubj+  h%h(K ��h*��R�(KKK��hR�CH      �?        �p=
�C�@              �?]���(<t@                      �?�t�bubhz�h{�h|�h}Nh~NhNh��h�j�M  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  (G?�������G?�xxxxxxG?�������Kt�j�+  �j�+  �g�j�+  j#N  j�+  j$N  j�+  j#N  j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  G�       j�9  G�       j�,  G@4      j�9  G@      j�9  G        ube�_legend_title_box��matplotlib.offsetbox��TextArea���)��}�(j�,  jw,  )��}�(hp�hqNhrNhshwhyj}M  )��}�(h�Kh�Kh�}�h�Kh�h�j  Nh�j  )��}�(h�}����M�j.N  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj   j  )��}�(h�}����M�j.N  sh�K h�h�j  Nj+  h%h(K ��h*��R�(KKK��hR�CH      �?                              �?                              �?�t�bubj+  Nubhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  K j�  K j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  G@(      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubhp�hqNhrNhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h���	_children�]�j,N  a�_offset�K K ���offset_transform�j1N  �_baseline_transform�j:N  �_multilinebaseline���_minimumdescent��ub�_custom_handler_map�N�	numpoints�K�markerscale�G?�      �shadow���columnspacing�G@       �scatterpoints�K�handleheight�G?�ffffff�	borderpad�G?ٙ������labelspacing�G?�      �handlelength�G@       �handletextpad�G?陙�����borderaxespad�G?�      �_ncol�K�_scatteryoffsets�h%h(K ��h*��R�(KK��hR�C      �?�t�b�_legend_box�j'N  �VPacker���)��}�(hp�hqNhrNhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��jYN  ]�(j*N  j'N  �HPacker���)��}�(hp�hqNhrNhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��jYN  ]�jwN  )��}�(hp�hqNhrNhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��jYN  ]�(j�N  )��}�(hp�hqNhrNhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��jYN  ]�(j'N  �DrawingArea���)��}�(hp�hqNhrNhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��jYN  ]�j�M  aj[N  j�,  hRC�p=
�C�@���R�j�,  hRC*\���hu@���R����width�G@4      �height�G@      �xdescent�G        �ydescent�G        �_clip_children��j]N  j�M  �dpi_transform�j�M  ubj)N  )��}�(j�,  jzM  hp�hqNhrNhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��jYN  ]�jzM  aj[N  j�,  hRC�p=
�#�@���R�j�,  hRC*\���hu@���R���j]N  j�M  j^N  j�M  j_N  �j`N  �ubej[N  j�,  hRC�p=
�C�@���R�j�,  hRC*\���hu@���R���j�N  Nj�N  N�sep�G@       �pad�K �mode��fixed��align�j�,  ubj�N  )��}�(hp�hqNhrNhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��jYN  ]�(j�N  )��}�(hp�hqNhrNhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��jYN  ]�j�M  aj[N  j�,  hRC�p=
�C�@���R�j�,  hRC]���(<t@���R���j�N  G@4      j�N  G@      j�N  G        j�N  G        j�N  �j]N  j
N  j�N  jN  ubj)N  )��}�(j�,  j�M  hp�hqNhrNhshwhyNhz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��jYN  ]�j�M  aj[N  j�,  hRC�p=
�#�@���R�j�,  hRC]���(<t@���R���j]N  j�M  j^N  j�M  j_N  �j`N  �ubej[N  j�,  hRC�p=
�C�@���R�j�,  hRC]���(<t@���R���j�N  Nj�N  Nj�N  G@       j�N  K j�N  j�N  j�N  j�,  ubej[N  j�,  hRC�p=
�C�@���R�j�,  hRC*\���hu@���R���j�N  Nj�N  Nj�N  G@      j�N  K j�N  j�N  j�N  j�,  ubaj[N  j�,  hRC�p=
�C�@���R�j�,  hRC*\���hu@���R���j�N  Nj�N  Nj�N  G@4      j�N  K j�N  j�N  j�N  j�,  ubej[N  h�jcM  �_findoffset���R�j�N  Nj�N  Nj�N  G@      j�N  G@      j�N  j�N  j�N  j�,  ub�isaxes���parent�hn�_loc_used_default���_mode�N�_bbox_to_anchor�N�legendPatch�jq9  �FancyBboxPatch���)��}�(hp�hqNhrhnhshwhyjeM  hz�h{�h|�h}G?陙����h~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh��h�Nh�h�h�h�]�]�����h��j�+  (G?陙����G?陙����G?陙����G?陙����t�j�+  �j�+  �0.8�j�+  jKO  j�+  jO9  j�+  (G?�      G?�      G?�      G?陙����t�j�+  K N��j�+  G?�333333j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�  j�,  hRC�p=
�#�@���R�j�  j�,  hRC]���(�s@���R�j�,  j�,  hRC�G��]@���R�j�9  j�,  hRC�����LD@���R��_bbox_transmuter�jq9  �BoxStyle.Round���)��}�(j�N  G        �rounding_size�G?ə�����ub�_mutation_scale�G@$      �_mutation_aspect�Kub�_legend_handle_box�j�N  �	_loc_real�K �
_draggable�Nubj�D  ]�(�matplotlib.collections��PathCollection���)��}�(hp�hqNhrhnhshwhyj�  )��}�(h�}�h�Kh�h�j  Nubhz�h{�h|�h}G?�      h~j�  hNh��h�j�M  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jfO  �remove���R�h�Nh�Nh�Nh�Nh�Nh�h�]�]�����h���_A�N�norm��matplotlib.colors��	Normalize���)��}�(�vmin�N�vmax�N�clip��j�,  j�,  )��ub�cmap�j~O  �LinearSegmentedColormap���)��}�(�
monochrome��hd�Greys��N�M �	_rgba_bad�j�+  �_rgba_under�N�
_rgba_over�N�_i_under�M �_i_over�M�_i_bad�M�_isinit���colorbar_extend���_segmentdata�}�(�red�h%h(K ��h*��R�(KK	K��hR�C�              �?      �?      �?�?�?      �?;;;;;;�?;;;;;;�?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?                �t�b�green�h%h(K ��h*��R�(KK	K��hR�C�              �?      �?      �?�?�?      �?;;;;;;�?;;;;;;�?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?                �t�b�blue�h%h(K ��h*��R�(KK	K��hR�C�              �?      �?      �?�?�?      �?;;;;;;�?;;;;;;�?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?                �t�b�alpha�h%h(K ��h*��R�(KK	K��hR�C�              �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?�t�bu�_gamma�G?�      �_global��ub�colorbar�N�callbacksSM�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ub�_update_dict�}��array��s�_us_linestyles�]�K N��aj",  ]�j�,  hRC        ���R�N��a�_us_lw�h%h(K ��h*��R�(KK��hR�C333333�?�t�b�_linewidths�j�O  �_face_is_mapped���_edge_is_mapped���_mapped_colors�Nj�+  j�9  j�+  h%h(K ��h*��R�(KKK��hR�C �?�������?TTTTTT�?      �?�t�b�_facecolors�h%h(K ��h*��R�(KKK��hR�C �?�������?TTTTTT�?      �?�t�bj�+  �face��_edgecolors��face��_antialiaseds�h%h(K ��h*��R�(KK��h/�b1�����R�(KhCNNNJ����J����K t�b�C�t�bjR,  G@      �_urls�]�Naj�+  N�_offset_position��screen�j�,  Kj�+  Nj�+  N�_offsets��numpy.ma.core��_mareconstruct���(j�O  �MaskedArray���h(K ��j�M  t�R�(KMK��hR�B�!  333333�?        ffffff@              �?        gfffff�?      �<�������?              �?        333333@        ������@        �������?        gfffff�?      �<      �?        �������?        333333@              �?        333333�?        333333@        ffffff@        gfffff�?      �<333333�?        333333�?              @        333333@              �?        333333�?        333333�?        ffffff@        333333@               @        333333@        333333@        ������@        �������?        gfffff�?      �<      �?              �?        �������?        gfffff�?      �<      �?        gfffff�?      �<333333�?              �?              �?        333333@              @        333333�?              �?        ffffff�?        ������@        333333�?        333333@               @        ffffff�?              �?        ffffff@              �?        gfffff�?      �<gfffff�?      �<333333@        333333�?        ������ @        gfffff�?      �<       @        gfffff�?      �<333333@        333333@              �?        ffffff�?        gfffff�?      �<333333�?        ffffff�?        ������@        333333@        gfffff�?      �<������@              �?              �?        333333�?              �?        �������?        ������@        333333�?        ������@        gfffff�?      �<ffffff�?        333333�?        gfffff�?      �<      �?              �?        ������@        ffffff�?        ffffff�?        ������@               @               @        333333@              �?              �?              �?        ������@        333333�?              �?        ffffff@        gfffff�?      �<      �?              �?        �������?        333333�?        333333@               @              �?              @        333333�?              �?        ffffff@        333333@        gfffff�?      �<ffffff@              �?               @               @        gfffff�?      �<      �?              �?        gfffff�?      �<       @        ������@        ffffff�?        333333@        333333@        ������@        333333�?              �?        ������@              �?        333333�?        ������@        gfffff�?      �<      �?        ������@        333333�?              �?              �?              �?        333333�?        ������@        333333@        333333@        333333@              @              @        ������@              �?        ������@        ������@        333333@        ffffff�?              @        333333�?        ������@              �?              �?        gfffff�?      �<ffffff�?        efffff�?      ��ffffff@        ffffff�?        ������@        333333�?        ������@        ������@        �������?        ������@               @        ffffff�?        333333�?              �?        ������@        ������@        ������@              �?        ������@              �?        ������@        gfffff�?      �<ffffff�?        ffffff@        333333�?        333333@        gfffff�?      �<      �?        333333@        333333@        ffffff�?        333333�?        gfffff�?      �<�������?        ������@        ������@        333333�?        ffffff�?        333333�?        ������@              �?        ������@        333333�?               @        333333@        ffffff�?        ffffff@        333333@        gfffff�?      �<333333�?        ffffff@        333333�?              @        333333�?        333333�?              �?               @              @        333333�?        gfffff�?      �<ffffff@        gfffff�?      �<333333@        ffffff�?        ������@        gfffff�?      �<333333�?        �������?        333333�?              �?        333333�?        efffff�?      ��ffffff�?              �?              @        ������@        ������@        gfffff�?      �<333333�?              �?        ffffff�?        gfffff�?      �<333333�?              �?        ffffff�?               @              @        333333@        ffffff�?        �������?        ffffff�?        gfffff�?      �<������@              �?        333333�?        333333�?               @        333333�?        ffffff@               @        ������ @        333333@        gfffff�?      �<������@               @        �������?        333333�?               @              @        ������@        gfffff�?      �<       @              �?              �?              �?        ffffff�?        333333@        �������?        gfffff�?      �<333333�?              �?              �?        �������?        333333�?        ffffff�?        ffffff@        ������@        ������@        333333@        gfffff�?      �<      �?              �?        333333�?        gfffff�?      �<333333�?        �������?        ������@              �?        �������?        333333�?              �?        �������?        �������?        ffffff@        �������?               @               @        333333�?        �������?        �������?              �?        gfffff�?      �<gfffff�?      �<      @        333333�?        333333�?              �?        ������@              �?              @        ffffff�?        ffffff�?        333333�?              �?        ffffff�?        333333@               @        333333@        333333�?        333333@        ffffff@        ffffff@        333333@        gfffff�?      �<      �?        ������@        333333�?        ������@        gfffff�?      �<333333�?        333333�?        ������@        333333@        �������?              �?        �������?        333333@              �?        ffffff@        ������@        333333�?        333333@              �?        ������@        333333@        �������?              �?        333333�?        333333�?        ffffff�?        �������?        ffffff@               @        333333�?        333333�?              �?        �������?        gfffff�?      �<      @              �?        333333�?              �?        ffffff�?        ������@        333333�?        333333�?        ffffff�?        gfffff�?      �<333333@        ������@        ������@        �������?        gfffff�?      �<       @               @        333333�?        gfffff�?      �<333333@        333333�?        ffffff�?              �?              �?        �������?        ffffff@        ffffff@        ������@              �?        gfffff�?      �<      @        ������@        ffffff@        ������@        ������@        gfffff�?      �<333333�?        333333�?        ffffff@        gfffff�?      �<333333�?              �?        ffffff�?        gfffff�?      �<333333@              @        ������@        ffffff@        333333�?        333333�?        gfffff�?      �<       @              �?        333333�?        �������?        gfffff�?      �<333333@        ffffff�?        ffffff@        �������?              �?        333333�?        ffffff�?              �?        333333@              @        333333�?        333333@        333333@               @        333333@        ������@        333333@              @        333333�?        ffffff�?        gfffff�?      �<       @              �?        ������@               @              �?        ������@        ffffff�?              �?        ffffff@              �?               @              �?        ffffff@              �?               @        333333�?        333333�?        gfffff�?      �<       @        ffffff�?        �������?        ffffff�?        333333�?        333333�?        ffffff@              �?        �������?        �������?        �������?        ������@        ������@              �?        ������@              �?        gfffff�?      �<������@               @        ������@        333333@        333333@        333333�?        ������@              �?        333333�?        ffffff�?        333333@        333333@        ffffff�?               @        ������@        �������?        333333@              �?               @        ffffff�?              �?               @        gfffff�?      �<      @        333333�?        333333�?        gfffff�?      �<333333�?        333333�?        gfffff�?      �<      �?        333333�?        333333@              �?        ffffff�?        ������@        333333@        333333@        ������@        333333@              �?        gfffff�?      �<333333�?               @              �?        ffffff@        333333�?        ������@        ffffff�?              @        333333@        ffffff�?              �?        gfffff�?      �<������@              �?        efffff�?      ��333333�?        �B8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �Nt�b�_offsetsNone���_uniform_offsets�N�_transOffset�j  �_paths�jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�B�                �rSl��?      ࿉��e��?���֠ܿ�;f���?�;f��ֿ���֠�?���e�п      �?rSl���      �?              �?rSl��?���֠�?���e��?�;f���?�;f���?���e��?���֠�?rSl��?      �?              �?rSl���      �?���e�п���֠�?�;f��ֿ�;f���?���֠ܿ���e��?      �rSl��?      �              �rSl������֠ܿ���e�п�;f��ֿ�;f��ֿ���e�п���֠ܿrSl���      �              �              ࿔t�bjm  h%h(K ��h*��R�(KK��h/�u1�����R�(KhCNNNJ����J����K t�b�CO�t�bjn  Kjo  G?�q�q��jp  �jq  �ub���_sizes�h%h(K ��h*��R�(KK��hR�C     �H@�t�b�_transforms�h%h(K ��h*��R�(KKKK��hR�CH      @                              @                              �?�t�bubjiO  )��}�(hp�hqNhrhnhshwhyj�  )��}�(h�}�h�Kh�h�j  Nubhz�h{�h|�h}G?�      h~jF  hNh��h�j�M  h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�h�jfO  �remove���R�h�Nh�Nh�Nh�Nh�Nh�h�]�]�����h��j|O  Nj}O  j�O  )��}�(j�O  Nj�O  Nj�O  �j�,  j�,  )��ubj�O  j�O  j�O  Nj�O  h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubj�O  }�j�O  �sj�O  ]�K N��aj",  ]�j�,  hRC        ���R�N��aj�O  h%h(K ��h*��R�(KK��hR�C333333�?�t�bj�O  jKP  j�O  �j�O  �j�O  Nj�+  j�9  j�+  h%h(K ��h*��R�(KKK��hR�C �������?xxxxxx�?�������?      �?�t�bj�O  h%h(K ��h*��R�(KKK��hR�C �������?xxxxxx�?�������?      �?�t�bj�+  �face�j�O  j�O  j�O  h%h(K ��h*��R�(KK��j�O  �j�O  t�bjR,  G@      j�O  ]�Naj�+  Nj�O  j�O  j�,  Kj�+  Nj�+  Nj�O  j�O  (j�O  h(j�O  j�M  t�R�(KK�K��hR�B�        �?������ɿ      @�������?       @        �������?              @�������?333333�?��������ffffff@033333�?      �?������ɿ      �?        333333�?              �?        333333�?              �?              �?        333333@        ffffff�?               @033333ӿgfffff�?      �<333333@        333333�?        333333@              �?        ffffff�?��������      �?�������?������@�������?gfffff�?      �<      �?        gfffff�?�������?gfffff�?��������������@        �������?��������gfffff�?      �<gfffff�?      �<333333@        ������@        �������?������ɿ333333@              �?�������?333333@��������ffffff�?               @              �?        333333�?        333333�?�������?�������?��������      �?������ɿ������@�������?ffffff@        ffffff@�������?������@833333�?333333@        333333�?�������?      �?�������?333333@��������333333�?�������?333333�?              @�������?      �?�������?333333�?�������?       @������ɿ������ @��������333333@              �?�������?������@�������?      @        333333@        ������@�������?ffffff@��������ffffff�?��������gfffff�?      �<      @�������?333333@        ������@�������?������@              �?������ɿ333333�?        gfffff�?      �<ffffff�?              �?������ɿ������@�������?      @�������?      �?�������?������@               @              @        ffffff�?        333333@�������?ffffff@��������efffff�?      ��333333�?               @������ɿffffff�?�������?ffffff@�������?333333�?�������?      �?        333333@        ffffff@�������?      �?        �������?��������333333@        �������?433333�?      �?        gfffff�?��������      @�������?�������?���������������?��������333333�?�������?333333@        �������?��������      �?�������?333333�?        ������@��������333333�?        ������@        333333@�������?      @���������������?        333333@�������?ffffff@        333333�?        333333@              �?�������?      �?        ffffff�?�������?������@        333333�?        gfffff�?      �<������@        ������@        333333�?              @�������?������@        333333@���������������?433333�?�������?��������ffffff�?���������B                                                                                                                                                                                                                                                                                  �Nt�bjP  �jP  NjP  j  jP  jc  )��}�(jf  h%h(K ��h*��R�(KKK��hR�B�                �rSl��?      ࿉��e��?���֠ܿ�;f���?�;f��ֿ���֠�?���e�п      �?rSl���      �?              �?rSl��?���֠�?���e��?�;f���?�;f���?���e��?���֠�?rSl��?      �?              �?rSl���      �?���e�п���֠�?�;f��ֿ�;f���?���֠ܿ���e��?      �rSl��?      �              �rSl������֠ܿ���e�п�;f��ֿ�;f��ֿ���e�п���֠ܿrSl���      �              �              ࿔t�bjm  jP  jn  Kjo  G?�q�q��jp  �jq  �ub��jP  h%h(K ��h*��R�(KK��hR�C     �H@�t�bjP  h%h(K ��h*��R�(KKKK��hR�CH      @                              @                              �?�t�bubej�D  ]�j&E  �j'E  jw,  )��}�(hp�hqNhrhnhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  G?�      j�  G?�      j�,  �)Residuals for DecisionTreeRegressor Model�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j6E  j�,  j�,  j�,  G@(      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  �center�j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  Nubj7E  jw,  )��}�(hp�hqNhrhnhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  G        j�  G?�      j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j6E  j�,  j�,  j�,  G@(      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  jr+  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  NubjFE  jw,  )��}�(hp�hqNhrhnhshwhyj�  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�  G?�      j�  G?�      j�,  h�j+,  j�,  j�,  j�,  )��}�(j�,  j�,  j�,  j�,  j�,  j�,  j�,  j6E  j�,  j�,  j�,  G@(      j�,  Nj�,  j�,  ubj�,  �j�,  �j�,  j�,  j�,  j{-  j�,  Nj�,  Nj�,  �j�,  Nj�,  Nj�,  G?�333333j�,  NubjUE  j�  jVE  js9  )��}�(hp�hqNhrNhshwhyj  hz�h{�h|�h}Nh~NhNh��h�h�h�Nh�Nh��h�Nh��h�h�)��}�(h�h�h�}�h�h�K ��R�h�Nh���ubh�Nh�Nh�Nh�Nh�Nh�h�h�h�]�]�����h��j�+  j�+  j�+  �j�+  j-  j�+  j�+  j�+  jO9  j�+  jcE  j�+  K N��j�+  G        j�+  j�+  j�+  G        j�+  Nj�+  �j�+  Nj�+  j,  j�+  j�+  j�9  G        j�9  G        j�,  G?�      j�9  G?�      j�9  G        ubjeE  �jfE  NjgE  NjhE  �jiE  N�_subplotspec��matplotlib.gridspec��SubplotSpec���)��}�(�	_gridspec�j�P  �GridSpec���)��}�(jr+  Nj�,  Nj{-  Nj�6  Nj�E  Nj�E  Nhshw�_nrows�K�_ncols�K�_row_height_ratios�]�Ka�_col_width_ratios�]�Ka�_layoutgrid�Nub�num1�K �_num2�K ubjjE  NjkE  ]�(h�hnejmE  NubjW+  Nj�,  N�color�Nj'E  N�colors�}�(�train_point�j�M  �
test_point�j$N  j96  j,,  u�hist���qqplot���_hax�hǌ_labels�]�(j�M  j�M  e�_colors�]�(j�M  j$N  e�alphas�}�(j�P  G?�      j�P  G?�      u�train_score_�j�,  hRC      �?���R��test_score_�j�,  hRCd�{L�9�?���R�ub.